��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����Y_��F��tw�p�^�=�����DW!of�.��"�"V�8��Ua}W#R�M�-Q�xq��ų�����#k_Q��?���B8I��c��l��{ͪNȽ�D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȦ�A�k��V��Af�{��b?��iY�c��Q[��|X@nl�Y�J:�H_0���k3��S��K��I?+�؋�}���b��y�m�i��h�,I�m=�?�C��/�o!�L��A�b$����q�]`���� ��ބZ|�[��Wq_^�ח�����̟~�b��-x�/��jRx�N�����A�s��cg�]�}�?d�� ^��b]}���͔�򐌹��	0�����>�r�k���Y��cd#N�N�W�>�ѽ�:�U�".8�> =x$i֒K�{��_^���Jt�]8X{�u�qA3���:���j�5�`�b���6w�5H+�����e�3(�Ꮝ')��r�1�b�=&�`_���f`9�MC�hM[��-9�B{�}\IG��O�Ҁ�żS�sZJ��� �*�����#��܋��D����9����g���e���놔���ʈ0��o����X1\�Sc��!(�HU������j�Ҏ�d�^�	%��������ϻ�U�J��/��*�vX0B�8.���H\%Vg�&���15?X*bXHV�����/�)����y�� z1o_�C����a�5�9�#N��N�]|��b��=$ǵ5��B0���1ɥ���7 ����B��h=]d���֢��]a���{��ɏσ�Z���PQ9!�̲��NAk1I�N�qU�<]�����J�L��������L�V�|�����ȓW���yp.z�WE�=;	���*%�[)��_�c��(�Q�:����h�j�"�q���m+��^@n5�ŵas|4��/��H�N&d�@a�������!a(�ٌf���^���5������7{�O5�b����]�-|��Q[� �|i9�@'9�F��^��Ʊ7��2�O1a�s��]Q�T���5̇y^V�Ah�g$�5�&�:� ��<���@��mzb@�rG�r���������Lg�D�V4�O~O"|��>���H�F��0�8�aI=�vJe�c��S\���E������<^"��M��ωIH��er�٣�E�@Ð����O�?�R��x�
}�c7ɽФ(�����G�ڬq�ۻ�a1χ�i�R�B�M�;Mn�?�S��vC���z�:�&���"�D��X��~�t��£�"��Ci%-=�F��K�h���/�k�2�%��u��Yp��UD�@�L,�ݸ*��߮����q�j��v��Ep�]F���1�X���H�'�c��R
)�ˣ&��+�tTgҲ�5�%ꟓ�;���'P��X~2l�0ٺ��G�WJ�;���͢o��v��׾�Q@D�=�Q)J
Ɣo�O�rv3�l�~+C�^˚�*���~�x(�7��㘿[��x�:�}�YM\?�*:����>��\
@�Z=�{>�	V�~dK�����<)�Ն�D�x��:�n}~��2�>{�-mW��2A���4�r}�cq�ժ�i��oˇ�G�GV�a�yӫ�R�u-�m/�p|_nU|����+h(g�o)�
D�cFl��;OA0`��<�@�ck�����ׯ��ZBFǕv+�L�Dʝ ZL���QcU��L��0�?ǰ�u����M#��<hzq`����S�0q�ȼ��5UKU͸�[\sB&$�9Un톒M��\���|�Kv���af�9�r|��+nw�ަ/=�X��9�-Vʟ;]֘z��D �5�Mj����Ԍ�d�֣sE8�s�{]���76�R�}�hc��RF�F��	��V@C(�9���#�u[�kPl�y1�0�}[��U���A"bj́��� G�N �ye��������t��J��RU� �7mH�Ԑ.������p�!#���kt	��[1&��������N��ks���<�K��bQ����I>�i�ފw��s0��1�|w=����+C&a���JR��o�`#���nƱ�*&3� ��*��5�K�����a�
e$?j�ș/��&�ȷw��v�$��E8LaF�NvA2��9W�?�)d���d)M�����xV�˲���s�Dm�0�*$g@�vdg��r�F��W�FS@�c�%Ï��tE����-�w��~�Lr$�g	Z6�-_�(�Z�2c�y�j�ҳ���R�R�$�o8>�.�x�'���SL���uR�9j�of2Z2�X��Ԙ�-qK�/��ү+8+S�y���PAZ��ZŲ�d��-����dh�=ͷ6�'
؞�(��j]AV�����������+R��ךejaޢ�Qz�6�4� s�kس�9����̱A���ޱ�^r����:܏lM�1i�lt��8,h����l�!�G9Yn;î>u�%D*���1)���+>�[s)ī�~��J2ɸ&�M�����b�?^��Q%8�;����i��1���ʃB�گ�0����8u������d�1��_��-��|İ#�#���8@]�wIP-Tua��#�z���`b9���\m(��4�����J�֌����nPadx��4
`��w�3 ����n��C�e����PlDME�����}�8�#8o�����Z�7*��Xԗ���Mb��QH�r����ʾ�(ˮZ�?��#ֱ�߬�� 8F������喔���
�F�+R���73�(s�1��cz�}�Ҧ�-�/�GV���8��\�*��p���>!p��Y����������Q;����A"_�pW�����wl�+=h��ӠS����hXgG���FH\�2�e[P�AV����v��]�k��хW��_�WuG��Z��O�N�W�J���q��v��h�D>>���aI���ob��'�A��l��*��*�����aI�Lmʥ����� �ٝ�ӧs�ʓ�}Q�Z5_��xy�d"�m{.i�������q����!�M:��.ҲY��S����E�;:Uw��MB�Z &��[�[�L�OLUj������d}+��4Uʯ
P'-�� ��+����,�xT@��S:�^��fO����So���PEs�a�8~�� KM3�-+El$�?n�o�J��P1+��Ӧ��~�+�m{�J�BWϑ���*yv�������"�N�JnM��\�!+f��|��v���oU^�-&�������Y���u�*+��p�^��(�:������{̀ΰ�KP-����8��$x�6�Sܱ��.��rF��x�h@3W&����Tk�� �݋�c��=��@謏���ȯB�.��
�<��$Y�qR��7،D�L��̨t���@�L�N*�	�P��v��C�x!2��'H璋�ex19j2"?4i���#���Dx�R^d���'�>�o��,I�e����˘U�~5Ds�j�M����d;�2�1_�'3��A���4����`���J�FR(�H�>F-;B�F�h~y��صI(14�.�cPK���}�D(n˂�[��A�6��`�򥴆��긇^�/8ċ�=ؿ�-���=�E�I��>]5����N��y�G�z���J�%FA|Q��Cl[��_|o�A��\��|���J${���usT�6]��^\3��^�7����0/7C��A�Yr5^��'�/�sԊ`�y_�|�9e�z�`�dD��J�rE� d�`�#�*J���%�y�f��D�j�@��2�5\۹�#`��L�E19T�_&�,ѳ�Sbi�:��
�J f��9��b���$	�V�r/�o^�v+��Ц=/B �������:G��q�� �A��6��t=b��\���=4m�<TJ1AzT�d�w`��Ej�{� ���f�m�����;�#O�dAc̄��&|6E��6�P�unϭ��Eu����M5�>FJ'��}���m�sLb�|V@㧽ڢ)���~��s��K�V��)	�6���\�[eљ�/-�6~��|],��x�O8� �)�҆��`m����懘`��/��,I$Ozþ��K��Z�^���S1�*���y����e7<5A9�uw��b�?�X
�iQu�}��|���z8?;`ZV#k�&��*����^u{�P�7�g$�l	)6W꾡�&2!η2x\v%�ϒ�i�!����x`�[��H�M�3����n蜗�L��Y���EZ�x<2�� +��� ��Gz/�$����Ps1d^�~��:m
_U��6���	��B�� �ز�dB�qU���|��*�is��yIM�Ğ�{"��܈o���`kK��<��&�ʖ��;�a���UIU*ӂ�\������S�c������!���`%;P�@o��'-���Q�"%ZPn ��ntc�vD��|�=>z��_���ޅ� Ș�)������s�����5�;������cv�F�KoXƦo_f掔">-S���Y�\1X�E� #�� N.�3W .�b�l�^.�|�>l�M{"jc2���
5%pB,_��S3r�;
W�n�Qz]� ��J0�(U|�yUrЏ�t"Bj�#@rp�*x�
�:C�~y_���/((�-��lZ���w� D�n"��
W+:p��1�QIf��}���.άXTREL�/��7��i� `��τf��͆��'���燑d�>�����.Scv�LX�����gN�Z�9L��bB��1��}��T�'V�����M�}���o�SAo*�VY���*qI�+Rzj�S25���`$A���on	7�k l>�	�	Rb-��j�𵽫�b�cZUH�|��y�T�)V5Q��&~l���J �c�dG����E�]�R�%ž�\�Pc��4
���u��{���Ƚ�[�� �3���B�-�R�K�ͻ8�=��T�(?��}0Yd�N�m���K�8��-�T��\�pS��f��|�I�-(�E�Bh�@i�a��� \�P#F��&;��ڔ&k��������g��K���ce���$����?�J�K�#��d��U'�ӱJ�)�&���wR����x%�2�:;�Oe&�z�]O��BKw���폾���)��R�z�z�q;�o0��E����t�SER�� ��>_�`���I�[��7��7�I�t�A1Ѯ���s0&��[) �jp���ا��?��ج$��$c�,ax;]*x<@��QQrW�����; $�D�T��ݷm'ܥ����$$��$�p/���M�����O �؏�B<�2xg���x>OL�ܔB�$�,j� H�T����Ū&a3{�۽�k�����\��-�|�-Fw�����3�J�2�]�``4��� Y�
�=v��p6�ˡ0�f��&6ҥ�����b�v�S��E:�j;oP��;.n2/v,������>X�)If����d7^w�]7B�A���d�����`��[��)X�����S0U.�E�X��U�
������8���]M ڈ��)�sA���R��q�`aCz����[�����/绠�PU1#@,�����Ю�]�z�oV�n�U��T^����|��X�����,>K�pShq���q��eB=�A����z����J�?l���ӌ)��د]�{L��d�8��OY�U[הkyr��߫ �,%=�s]��Q\�pZrz}����^�4�r�v�
�~�X���������m����Ӫ�{eS����_����u�h��4d��͚�v?��cs2$���+i��\�FM�r���*k�,��[��U�0������@N�������#���Ɏ�WXAo���Ҋ�l@�9'��U[�\#�;�Z�8���oY&����'E�D�n/TG]�0�O(g�\:��J�7�"ç��\ %��as�y��*X��iE}���^X�d���l'� q�<���m��D�Vl6!bԨ����me>�E!��h��d��O[ų`�xiUIjl �?�5��,��:�Vɞ��j�P���h**�H��0��Ə Ԛ���ŗ�= ��[[��!}n���}ߔZ{$hݭ��}M`	�q���语�/�p���aI��Q��	?x^A����حT��V$�?�����2=�$x_�+j:��xx�E73�Bt�|�^.I��B/�l�>�F�����Q:�vT�c}���*v�7���rT����ʲ9�i��W��3�Zn꣝�����>�Dq�P���Y&_0��fϠ?�):�<���	j4mL���9��Z��-��S<��nZ�W\=_5�����Cs,����1U�e�z����5�x�9醬۶�Ϧ���9����#��(�q���0#s����~����9�0 랑;sK'R+`�!��6'F|1�SI��I0!1�@�Ug�Q��Qڒ9�v	cH�W!RN��6~�~ ���z���*Pa>��Fū83򿽭��Z���{����U��§-�ק�Q.��ҧ�g*�󬰜�n�1��A�5���|<�L�H�w���]���z�5V��JL��o��(dN��h{+e9s๠�^��O�5�eM���_\<7�{[��rBf�� ]��J��K,)�y:F����j't	�[=F���0��߱[Gā&K�I��I={���#�-2'�=H����̈�DO�x���e���Ǩq��0d``'Z�{�i�tVǃ
ȩI�}>�ʐ��5H�b~�2��.n���Y�w%J��P�H���1����˴K������r1�Z��7ƭV�@'���6�:(�&�0�#�0|���I����B[+!\!��>L u���i��p�^�����=�k�\MN�|�W�' ��0E�ƺr�ڭR5Ķ���y�;6�玊3Yg���@���\ ���e,�����M���!"�|��~f�h��,=�S6G�E�2f&��T?1�0��#P	]�_�1��)�,�g�;`?��~�#j�T��؋���
����-�vv՚\�]��7]��#$x��I�v����#N��Yg�H.��i^�lƥ�l�<�(���!;��H؍9�{�W��U�b;,��ft� ���b�?v޽�"QC��ڻ�o0���;��+��iZnr����EJ[-k%"��7j�l�.J	�/ȧ�@�f�;��&��YMjt'�w<:�#���`�7��ܨ�aGl���SEO��hKF#?��A)�؝l ����C�H�IY��ֳn�����JͿ��g`Z5�g-����S���7�E���r��pÁD�� =ry#��ɔ�X����_T�e�x�G%
��k�4oػi�N�t���AN�������alHh�Ԫh��/�}�҄@���}f��.��J�X~�O�������E�N��i�K�3�/ÜSxVL��X�<���I_��C��,�(��6!�����ɷdTV���,/�
H��~&�4B�T�>q)�V��0��6�8؝CC�\�)�
%-9����B����mL�o�!6����Y�B[eӸ������I��C�����]�M?��{O��zdӠ���5��WZ��l,w3[�h��OE�*��:՘s1�71cq�ڡ���NX�4�~k�`��kU��d���Zx��<���o����\����άs#��}_!�9NT��,g��ú�rm�V{Sx�����g{�U���O�s��ʲX�Io۩ʅ�)-�]����^�&�*�F�J�6�i����J��|0	jL�C���Ӌ�1Lԭ]j�';[���;%O���`/c�yA�j��-����K�;�+EX�O�'q�iǢsZ,RB{u���U�6��}��O�7�Ў���`Sq�g�q�[*HUه�����$����z2�U@#R%ɬ�>�l��g!�W��0�9bcnn_���[ωKmd,�BlI�K���Z�h���m�7���w����va��X5�I�c͊��9Y-�OMy��J.k���>P�; �a'3Z�p�QX@�jJ�R�ch�N���W����
��}1�烼RЋ��7M'��Z��p�*������V�J��� �h����B��ǚ�m�x��{��nc퐄A�+f�QK��vt{�sjUb(;=�0 PR�
<�m�e���\rh�a�G��/�A?�h;�1�K\
Q���m��o��4��P�;��~������tW��<s���\ls�/g�]���6�c��@��Mx;����#)�gKB���܎>������d]=��,���	�&E@C ����δ`�?!1h�.RYXWU��}V�z��KS0��.K��� D��Ŷ���#����<�!��Am)�I-El��+�jdзIK��Z�k�Ն�t�Q��ޏ�VC���0�u��Xɯw�>�zM'EWB9����5�;�2`,����������x��������G|�T~����k`�p��mQ�v�֯#5*�M������y9(d+ؘr�mb��^v�ٍCC��6{����&0`����i�����N[�U�qÄxac<~�W"�NQFf���\]�H��