��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��RKj���B�}Φ#�Q�%���L+��*|A`Bow�g)۰a��Ԇ�Tv��k#�fU���yx#2<s�����_I3"�ꕳE�5����jVcE�����"*�k���6�&]�ƺI,���!�s��S*��y�v)���lA�$���/�����V3�'|^1]�t��4��6�y�я�jx����؄:�&�C��2h �C�Š��{�)4��Yz�]�u�eW�թڲ��QM�YSÉK��a�%�.�q�������B�#�u�p��仏�� �I�.�3g�g�$���Έ�?-vx�T89�Bp�������/JCNJ�xf�Op?�9��C��:�]4;�����~��+��9#(���$�>V�oH���60FuM".���)x\�5F��ͷǛ��=�k�S��?���\Wը=7C~�s�X��k��R�b:�/���][35wLmO䧭�Pj�K�Ⱥ��t@U �Ō?['��z�	����BS�4��d�P�+�CW�(T��{]hԖ�����%�3������j!?�8��ى�͑zf܁�E��N�0_J��f�_��4��"��~�jg��:x����LL@���1ȓ,��Y���S����$pԆ�&��9�Op����%k+��JgY�u`��1�2@!��5C0j�$��&�T��l��wm9�R�G#n�����Ol��vݜ�	c�7\g8��Ad�S[J�x�hO[ D�"��h�B���d�sb6
�=�K�~���5Lv,x�T<5��d�no�R�`ϔ/r��g��1`�����)x�uI&,���ؽ�A�ҝ�B/�TF���w�;!���*��z5)a��Q&H"om�]�1gSi���\a���6��b�`�ɉ:�>{��4!1S�ܻ��I�V�Еj��d��E.�`��P�����	��Ͷc=���YY;;�d�]�dw���q�����s�hFk}��q�کJ���&�N��@�&ܿ�ܰ;�R�>.n����2�u�d��	"�Z�������l|zE�{���8>GBrnJ���1PJ�^Ғ'L7m�,�j��G+����^fv��,xNQ��":������0#�M\җG/�lT�'|�e�q�$�cGA��b�Z	��	�Nq88L
ٻ�
�V��T����חB�fQ�3 �
��Cv�[� ]D��3�\LV"Q\����z��:��Q] ĕ�/��M��rf�:q��م��(�8�5ר��κY��BO��O�4ޥl�w)(��_�a`��H��f����p���"u���n��p���6����׳�~�>N%��;���
v�����h��!�C�/��5�P�n�D��5,���0u���^>�u:�q�*=�r�7�/G�e	��y@�f��M��aݞ���X�O9W�	��	GD��$�fD�.H�j�9��HZ٢<[(S\%G�>ꆌ��rnʷ�U�[.�F�Q���|����?5�-E��R�����Z��`+]sB2x	�.�j�s?��������9}�?�M4�'7р��T�oUL�h���t�g�T�l��l��5��O?&��A�Z�X��쥕S��oS$����x߇��Z"r�>���Gc$g&���d6_��g�3��L?�a�����paPP3h������d�٤����*����(�i�
V'�	��t�Q��گB����ؿ���+�gH�G���F��$yv�]���=�[��)���!А���[F�{�csɋRE���&|z�kx�/;Z�%��6=\���6TX<��#f��C�I�ȍ�FMg�,+'z)��E��:R�z��o����J���8/��o'8"h����[�^��Rҿ� �[��`��-�ﭏӝ<_i^{�%HC2��T��&�I� ��aLF�J~��I������C�
R�Bq������2�pd1 �v�;�����/�ߥE��	0Sfx�Q�Ϟ����2�
��Y� u`��x>T�'�PJ�є�&�4�zBgW�0�P��>L���*�G�)��X"��N��]�7��YM��\v��!�MH�':��Y��J�r�y��.�6�E�F�)���C������!���~��Đi}��>�Y�W��M5�.t�
|t�����?g��D����G��p�L)-'�Z��q`�f��UK!�&�ć�f�� ����\��i����DMu� O�L�9���0�R�CT��m�����M�f����[��(wE>�"'� ��m�Hy.%��h6��q����F,{b��	L�J�]L�a�QA}��;�mT�q�h���D��RBb�U)��'"U����Ɇn�Ϡ�B:1��m;Eߢo6�j7[����GX��"��v�_��!ʃ�>�|tc���w�+DC���<,�������XR#����F���ޮ��S+c�Q�my�������t�v���Ϲ��s�$��8�]�|�����v0F��\~J�;�ݾ)��"#꫖�*G�˴�O�*�wP��n���ĴlQ84���LȾ��W���M4L����Wf���Q���_Y�ő�����-v�'^�{$a/��{�N��4]l���w��5~v��@�u��L�Ԅ�ä�!�`�q$ �	��dUH���ʉm�*3r���?D��g:X�epkI���cü V��;��>s�8�v��+ׯ$\۬��&�� ��_�c�,p'H���m��!��y
������;�{2�֜8R0�u�� .���M���CUp����_�\\�$0j���K^����y�fq�f���v%����E���4��Uu��Å �%�ی���H�(�ճL��oT]]�L(�{˯�+�{�
�݋]DL\�P S��s��jY��,bh��@���DzѪ(��.��A��~a�-~q]!�b�,0ɼ�"7�±i�D����YFBLSB�&�5؜�#Ԗ��- L"�M~Ǭex��U��� �CB֞"�<s�(c���A���>�!�[�T0���k�� H�)���������E��Z1i��5=�=K�ӳ���r(��oY\�r����k�,�S��9�����:/H�$�@U���`	.Q:57gO?��"��
�
|�P>�,�w8�F�!�;k�z|E�.����&�ݳ�@��)�~�ˌ��v�5a��t 	��,D@��9���E�xM���x�;}�rC�cL�q�Ovi���b,Ѣx��BWD�P�9�v_�$�<!t�pUSjÔ��ZdB<�y��.2RDP�a�0#B��\�Rq!2Z��NQ�HL�C�Ws����`eP��gي�f ƨ���,n���`�[y�o���?s��T����{������|O�5��|�(9�b6N~4T:��E�u�����QcS:���.:��;��bXSp8B��Ys+5�E!Op��[��¡+ɤ<xup �]G�4��+P?'�h��|�$�j�FB����4
��1P6-o�=��`4��AϏ�r+���@kƺ�[)�$ yLv�ֺ$�����UE5��%��� �ul_�ёB��jpd��Yj)0W�(rO��/y{���[0چ��Ŭƅj���@�=�2�����S=9���Y��H4�3S���LR"���&g��q!�ؙ��E��
�®\9jhD���F�ڭ��dF�5�bLPU�z#���*��w��� �����9��'�1ßJ �3�S�%��:�e/�Nb4ў9���JE���ض��2����R��+ߣͧ�B�ٜ�(st�`pk����⃵�V���	���"�ݰ�C 	��mZld(��P�m0���/m���(U^��wI�F'L�@�$3Z��d��[�����ֈc^T�XRds�	� �W�B7#�OhN��@�Y� ���K~[A�j�,�q�i�9����^Zc�\T��fJ8oL������l"��_�8B@nQ��Ŝup|�X�׺bN��o�!~�w��W����R"�5q��G��%��n]�ft��V6C��*����@�|�$�:C��T�6|<�|���u\{�Q�3 �XQ�����t�U��Php��ܣD�� �gj������HB?�N��AS�J�4>�;)�"�H
�5�����zjvK�c�+�	M���= �+\�0�܇���>,�_i�{]��D�\�Mꯠ�0�n�&H�|gEY�ҹ�[��clT��s&�E�M�����	�Z�P����4�ب 	;�O�-*rK�3U�F���i�%%��\�
���Glq�;ӡ��`8d���N"��u�`�v����Y<�[������g�f�*�����j��X���z�
h�O9�ĬB�;���/L����,�'_�h���?�)�U����d�,)S�+��cp�Z�/��u�4W1{G�<R�6�g�Czv�R|2tc��sɭ����nN�`_��(f$����}��|�`��I��mn�M����P�Z�ek�]-��<�E��O>*+A4�iAu�,'v��`�m\;�i9z)����u��F%L�E|�U[�������u�}�sDѕ�?��"�s��*�3����1��Q�{���%H���.9���!P��C�	�v���a<C��]�q3�SCԑ�T
2�����4�B'�������U&��OyU��n� 8�y�I���@�dv��}����l�-(<Z�z���著���ckٛ^��:D1���J"��$$�`|DsJ��x�-��͝s�]����J�V8A�}�Syx�H���~�g�L�+��B&�H��}4��I�rT\J�Z'���(� Mi�Z<	�Bv�C��1���N�ڌd��3l�����:9�4����=��k:�F��ys�Ԙd5�!��Fp�G�k���O�טq�-ܜc����G�&�����`Oݨ%�ѾتR����RK�,�)`pʽXb��zCc�6��\dN�)��w��fK�W�M �kT��v�|�����ƅ[�/Njà�Kw�O.�V��ݯ��{��!�<�!<��T�5�5
E�گ9G��Pu��C���7� Lm��+3��\1$�1��d���gi�۷HE�P�)���SB��T<���%��%���NY�ƥh7�ͦ�To��g\Q"R\6��5��P���Ɩ`i���-=��2��3\g�\q�Hz�͐⨒]�iN�q`:Jx�`Tm4�-�f/xB�9l�:xR_�Q�9����G>=�w-��C�����ŉ����"���pY�ψl'B�Av�ͩ-j�m�%���0Bv������b ��@gk,�� �(��&#��F��I���9�M����J���Lۍ��gķ�P�ӳ`��)�K���#�5)V�U6?$�!������]7N� ����.g�.�?>t��&H��b�O���K>�lzn������8ҺϬ�{�<p:��az}���ۤ�J�*>Y��*��e$��u������W�;�-���=U{�VN�IK弅�^��P��R�#�C$��		���l�#g� }ϟ�=>qawsO�7��b�'`��(J�
���A���4HPg��B��DZ1����C7��v"�N����+��7�)��c�¦���#��eS�6h�5O�w�A8��b*�E=�du�^J�c`5���V$ϭ�=	�uɢ�*X����������1��kP�1�7�:�,�#��~��D7I������`V�z�L�HH.,B	�P��:��6ri��^��-�� mm5��I����Yx��'/�G��C��_ě�v%��8+e,d�t��c��������A��V�F�l�.�L���&��hW\a���O��߻�w�WG������6W�U>��i�1$�8��.c��1C�˼��'(`ĪZXv5��@� �
������/�3e�1nza�8��j+��Nc���d�=n���� E�('ƪa�wm`H� �	�b�n�La��7's�W�ױ"4le]|h��%���mx4t���vko���S��[����b�ח��ܝ9z�"�qU����f�M��O���	�����K���$(�o��۸���+��L ��L���\ɒ�h���7�rU�g3?lێ�K��W=l;Fo�Y�ycy@_�U��u��Z�����?q@�E�a��7w��6��/ />:A<�,R���2��U4c�l�<��ZK�"�{�?�:ɵ�_��&pߢOU���
���$�`��s
���ԧ`ζvx󶓸5�M�a� �Dܥs�Xb����ů9�/��;O����jx%��G����m�y�M�bß�W� KM'e�l��G���?��[�]�[��yR��N�B��a~kk¬�X �����F�V$�X�Y��@���#�rj���SV��ٮ�l���ƹ�_)�曃�����y�U	�r+�:x\�Q���1g`\ꄝN�?!H&#�&��ĝZ+6���gR��$|��'�/;g��6�����%�D	�����>>�a�-"��-���K)�`��kgM���!��iO޹��F`<=��O��j�7�"J�qj�M�:E������C�IVs���inNh^W�o0�΅�ew$��]���mx�D��$>�m>��VEN&`Wa�-c� 5A�&�!L���0��d�Z�i���հ�%��u��߈��7L�`����"\������ϛ��C��h^����~l�{>�ap�1VSO���A��<�����y�8J�e�ޤ�+ c�����-��f�P�������[�H#��4��f��PQ���n�%��5��r ��9}�ْ��a�������^��	���걋���I��ǅ������3A��A{��f0|3�P���x���"/ݤh���|���ȏG7�;�EW���>z&6�ӿ���A�~0.	�r5"$|��nc��3����O��E����׍2���l�k�'/I�Y�r�*�H���CB�p�c�} �/G4���i���;d)g�Ζ�ֺI�$
�*F7��i��_Q�_:��S���m�.ˊi���5��{w�Ά�W���.]�u�
�����<�Z�W펶�L^���3���Hڎa�!����T�^��o�PC2�co*�`ާ���V�lۆەQ�Dn7�����E���0&�����r%Z�ӡ�I�	^P!�f+�!'pT�)�Pe�5�H_k�`=���2Տs
O��<ϥz��f�q���c�x+��[D*Y�_�s)j2
X�)�If
�HI!Ԙ^�2�l <�R�m�M���xh�6ʮOӋ/��E���$�U_�~s|,h�1�A{Q+}N�9�o|�����A��r-�?�쩩3�)�#�(�R�O�/Ͷ@���K��N �	�gS|>s����&#v.�gZ�r��NB:��ђ=��[f��m��mj��V���M�XG�
N��g�W���?���_��ܮx�*v�f3���tJ����iA�,4���M��d=L��Yb����eT
��;JB���r+Q�����l��+��q�i=��Z�mT�EC*W�?jE߭^H��G�I�1��?�������	�.I�l3WM�V��i�0��z�'�j�����u�ت�J�ɖ,[j���P.s�W��?���٫.�d}����p��ev�xA���*��������0�Ɵ�Gs\���?Y��jq�B���>oLGT�q:U[��c�Q��!����5s5���+-K��SO�3��1���4���*��e��I���u��$�7�q�i� գ��p���!�:����~@�L/���(�����"R	�dѭA�KG�'.F����2v�#�:����1���b��/?c�RZ�WYqǸ[6Jݵ7,�����k"V���
� �IK�U�!�s�i����67�k��e��g�ؓ�K�a<�
��{ (_���J��f�j�_c4�{��3�jO 0�片:J-`j�˱�޺�_�����u0@H�S7�wCM�x����ɚ� �/
ݲ���F,�[D��
�N������J��<���V~:Ǖ�)��3�e�����5���7��ݮ�t~���os�۬%�~����P)ED�&�q�V�)hhc2~b��KTh�)��0�G?"��VY�x�ho����~�	����(]]��bH:H�z^������$�oYA����S�Շ��@�N/cX�b�b�?m�ŵf��Wl�6X��4�۵3ƕ�z���
����J���os�)�E6}�X {�V��#�"đ�oC+����1*F�����Z�10ͅ˺ga33u�6b�D~W�';���*��^���;=�@ԷF`܈Rd����?:\3�!��v�+��35���#|���Y�1�^c�H��i=�,�7c�����*"�^<Bг����gF
��0�Sp����N�@gF�oN�
�w��LX< �l���8a�X�Ck��V�X广�M�laTq}�j�9�ɵ�Q!G܍:I��7�*f��0U�>am���҇1�:�]�঩���㻸
�`�|�d���l��{8�!C~z�ߩ#=��V�ߡ������ g�Yb$�\�(��Ҍ�8�[��̇A���nDK���ꚑ���*�I�Q
�3���V3��vqTy�L���b�A�٤`��ңN۠u�z9������^��A�̩K�"���-��NC<_��<�D �dj�~���Y\�]��K����|�ym^��\ƹGE����Ԝ���Jĳ�����Y#s9�'��I����VSxоE�RZ��
B�o�s�e��je̘��*��]Mz�E��$���4ʰ�#�?�Nq�	#�-���}��J&x.0=��@5�~�����A#�u�X��h8�;ՓX.�H{��Zt�ZHi�zN׬��N\e2[��i$Wc���|��RG6�+;	�L�ByR�`%W�K��0����\R��TV���u�F׆� ������']�T��%�l��D-������Q�H�y�����dԹ�h�ހ��J|�z�-=.du��� ј�NP�^N�eĤ���V6�h�n�g(��/	剀^��@�8�l��j�<���]G-�:0�E&� ]ܜ$
ZO��ܖ�4�1�9�v+�ߺ�W���܀DK�JصvC�
����������E{&k��>�O43�N���(&I�M���nR�V��|䷆V16�7>& �2�u�?�mR�DpBgJ���3�>oU�[����O&�ua���	�뜃��qZ�$�{#/m�B2�MK{J��e�>kܧ|;}�K^�%�B�Sg�/[������80�;kd Mc�C�4[c�-N��5Z�RfM�f��͠В��q��p4\W8��Y�i���:{/�����Q�Lj�)�&,Z-�����R��l�8�8�O����~o+!���+!F#��<-��'v�tf)�Q���*+�H���9������۷T9�'�ʐ��HF�&�xyƁFc��j��q�l�����A?�2ufm�p���1`�b���	���4Ci�$d$[���T��:�e���)��:;�	F.{�ȕ�̜g���\����b9�Z�k������b�;�wB���u�+�"Se�����Q_�L���M�K��xmM�̫�Α�M��	�|4�%$��g�kf9sUt��F"�#����ƚ�;"�3bRq5�wY����l<��u����,7K�h�b-����vׯ�}%����D�_�G�\�y��m�9�t���#�k?��T!FԨ߼����{$ݡ-Űҳ'�������0��љ'�0�P��TO�ĻB��i'K�f��Qt*4`!	��XJ<�8֚���O�-�4�/��+?W@�1J�O�V�	�IF��<z������w��ј���}Jk ���:i��X'�'�����^%R��̧k�$#�:M|�U�l.��P��m���=S5!���^=E1o��%A�-cH��CZ�x��q�N,��a�I��v����#ʃ��;�VO\���	SՈ�M&H�"���6i:� ����IƳ�e�VL~�w�Q�Ъ{���l����$�.��n1i�骨�`�Wң�g�[T3$���
^F	�v%~�j޺��`bi�w4��ʚ�U�US�D�$�<����e�{��0��[�nr���][�M�i8�f�s������@x�"ɋ�� �]�gph.Y�Y��(��Tuk �	�Չ��?�Y6h�̻������=��	x�-����1-*)�>�����.'���j'3AS�;�؁�M���h�nֿ��S��]r��T�Z�7kF�Xo�h��WΡO�༧���_0�S�è��Z!ɇ:��%����z�B0y�;�Lf���q�Z	��������[�:���![�a���*���[A�5��#K@:2�:����t�	5&
�x ;��L�=r03����!�5��m�zG8���>��aK7 ����(�ٕF��1}�<��~Z��������![�Ӈ�5�f�E�*�����R��/��l0���ƃr���r�c��?�����N�7�������� C�r��7�f�����&����I?�A�8	����Ѧ%�\Lb!��ΜZ���NCD�A���2��;��)t�72k�LNjcݸQj���Y�E����a��[h���|"tR�A�h�M�ʑ��xu�,�_W��)�NQ�X:|ffa�b��ixL�k\-x��N�tr�*����Eи̛���]�E1��a�ܤbaF���R]�fuPJ�F�s��%��%�}���?qՂ�g)x^�v���f����c�D!k��&坴~�K=��)<��_�j�o��V�$�m��U�;>Q�v��w���eb�==��*��+W��S_�:���A�"�F��YzP�
X�U`3�-�D����X!g"��hcI%fo��$���jp�҇S��EtcM*ބ��ɣ��a����	�[D��ȋ�0��K�TAa��o��<���Z5���:�����}����>!�����zS}:&���>5��xV�������m1C�-�,%��O��7��VB������}I���Cʶ��k��
	��Y�������#��3\�8��į�S�Rb��|:0ZR����?�<E��r��v�)/ei�k\"_��pHm��]����#HA#`0��[f�V_��?����x�y�x��I��-;ë��ɥT �槂����>�\h�u]���W�z{T��ա�b�-���{�#��]�6�E�e,��0U\m������X�z���Ym`^�_�ա�ph��1@�WmՔ�d윹�����y۱n�r�8M�I��c�=��\�i���Pw~�
k=�#��e6�kp,�I��oNv���VW�Z�������a�[�K���kr	R�̬�^i3�H*��D�Ҝ?�u���<��n��r��)������[!���E3�n�4� ��+��Ơ�..%	���դ�s���C���X�<�ӏ�PAĒ!��x� �^�7�C/.�l	���o(�1g?e��j��p��M`�WxSgb����)�}�/��l/3��aH��}��a�8���U�Py"��t���&>��;��s�{h�YXa�"ѐb��"�����M��N����(���n$�b\-J��ŧ�JV���o��8�H�.rG�����'ͦ�
㻸:�kR���>�����_�DN��R���\��A��B�K�߿��ͮ���Z4I@�سޯ6?���ݷ.~���o�J�舻GK2�=G�wKt
�6�4v��hoڟ�z~r�����=��>�#i�Kݮ|؛�Ŋ*_������9�:7����w
)����%W�����	�e�ڻ����
=��]�_NŸڻ+H�Q�N�t���J.�.,wg�m��*ߍ��X!�-*k!�z��r��HA?����'5�2=c�<��A8�ߪH��)�z�i�j�噾�!�e���{�f.�J�,P�}?��C�[Q����R6����P=/��MU�^vUn2��v��uOp&��-f�|��ƃ��.���dsy\si?�g���������;��#]����D����\$~��g__	�ȷ��A�/�,B�[�<����}{}���y
G#}�[�֭yipy>�M٥�Fi�F�4ps���a&�TW���<��an�"Y��H��Ǡ��y� |H��%���I�)Pе֤��0y%0��W![*ͻv�8bHq���^u���#�x:ޖ";P'Gvyq\���5��M�ȟ�Z�{��Ֆ�"��R㙁���:s��(�GF�kNo��J�&)�-:.��QOg�E2n��B-�u�Iĸ/�f3��$�p���o!~�z���u���Y׭�/��A<�pdL�\��J���(E����f(w_���w�D�dmL���6���Sz�4��g<��|m�!���2��a�&��ӹŌ�����\Q�ՠ��(T �s�'�H]K�W[+�軝����l���J>���8�����4�̵/�G��z�pPq6%�J�c�hOk��	i��/M
O���R��Y�n/G׃u�T���֟q�n%B��u�H�4�?&�#��rZvh�>�%����i��� ���)�'=~�N3�����fZ�]���$�g�ӕ��!��ր �W�)��/#�N�D��ά(h�?��䑘w�r���gYEI	��L=�^Fw�Cl���5]�d�{R/V�P2�{�vA���R�{�;�r���gm�#���S@��}����.�ꉣ�9D�w���Th̠�|"On�L� Ӌ�ل���|�|��c��X��lI�!C�wԡ�'neJ�4nn����H"C�y��beOV�mĳ��Ҷ0�������=�b9�~ˢx��v1QP��H��*�]j�ǣ��(5o]�\�ܹ��ڀ�Ps&��C*plK?h�	�.KЦU����t"������2qeQg��ml��\��c�x }���9�oV]��t·Bo��m� �*�~[�o��	�!m��F�䭻
G6 ğ�S|� ���wN��Ƚ����1t#=g'�	��F�_�s-��y�P�:�s(���b��EDg�W�{wJ�KO��t�(��H*�%dǲ�ea�P� $�u�R�\�N�;��c�f��{�t�=���uՌ_\�0#�e�Iڠ8C�*��-�g�S���wC��Q,K��-q���W���O�0f�]�:h�I��}��t��_�ɜ����B
���ȨةԖx�M����kX�gw3��e�v�ɿW!��LÀ�qIAM%p�xP�	,;��v8Un?�j\R;;ȯ���zJ�
�^U;Ly�l8�<���JY` �6�ZTYlM�?@5V'=K?+C�mb�;��	�i��"_�I�Y�UZ}��^Z��jb�4���1GώJNo��X��v�w�=�}�ϻ�rk5u!,	G`�淁��0p�����������1� K�&J�M�&	�}=�Q��^v��P��r`��"��G��onA1ԣ�=�N����ܣ��~�������@���^��B*����*���d�I��}��x�*u+bb�U1e�)��?��̭��YM2�i��աP����pۛ��U��bJBM?�0��,A �X�T�DPN��������TD�����g���,-W��(\k���v����	��9�y�h�x#\Y������dj�Tk}6�DL!�4���e�����Z����m�qtM]s�&�,/��#���u�[`��'3\��6�}�ų$p���)ǂ�w�X#	=���8W�N�ֱ���/I�@��M��U:�94����f"�
����VT�Ʃf%��"�uAk����u�C?�ص�|2}X�a\�o���R���%�s�w��b�ț"S��u��{Ӂ�hp�Ça6��|O��\ݴXW��`�+I�Y@f��[y�%*S0��=�o��p�K� ����[������>ߠ�{%�w�K G� Mz4b ���n"(�`���F�k:��a�������