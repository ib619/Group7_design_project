��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]��J�/�f�m�G\�t��Ʌ?-*�хK/��y"\1� 2���I�M����Ӆ8���ph�;%��q��g`��o��4bs-�����Χ��1��Lŏ�_�����#*�t�p�𗚻!��!������{,� @��H�X�4���;�ʻ�A��o�kd�'�;��K���I��_F����x���l��'Au���
�M�X#�_6	��G"��
#&Ç���!����Z��v	���ļUr��C�����p�<&�i�d�K ͏��wG����8 ��ȯ��c;�٢Db1��$�5D��JTK��k�Lc������V�5�T�Ф�1��۴�g2��#����L��Ƈ+zkoud�b�7��"?���[�,�=���� ���R��\l�K�r�M���4v������:�K	!�#`�e.��VT�W�qn����.��K7w!�uJ7����~T�>TLc4�	������X���%0����a� ���bE�&[i# D늬�$F�nJ���L��@���bu09{ie��䯈~|���{���+�ʎ�H]?��Q%18���|r�1��lؼ;y��;��� ����J��RKo(O}ޙ='Ya� ׅ_el>�Oq�EN �����sJ�VF��L�^XՆD��=�pR��wd����Cۧ��FWl����-�B
�\�����g�j�I���6�ap���ȋ+�}�%��'�O<��0�������	R����6Hb��s���
���.!��~��Q���]5�15�^��L~v�jċ��HA��z�1��U��2i|�<�e��Z8I�J|��� ����K�x]����%؜�LB�d�A^'*�!5�K�<�E1?�i�V�\0��`��ǹ� V������dw&o��i�'��W$�MY�<��l�f�����RF5vSMm��ށ��E� W��j������LG?��4m��kd,��_��5"I��B55=&G�W׸�١�Yx�P9��@�#�P��$���C��s��q�����w��@����d��F�?�a.��	^W�WT�߄9 �U[�)(;Q�A�;-�;���c0�����3Ogy��ڶEϾ�����-YPn��D�̥�hk����l����3�\�4���KXP�<d�����e�ܺ`�����;��k�j���n�/S�� Z���I¿�5�|��Y���S	
��l1��Sc�:�Q��!�T^�6"r'6&8�J�z�����"��TVD!��/.�Pĳ0�c}α���ǖ�[�d�#�E$E.0އy*��j�ib���U��V*C`v���P=�������$�XEHHPi��D�����;G1�H��^�,ގ?(�˧�F�O�fWQpzUp�T�-Ump�f��zf�n#��������M�|)���R��K�A�t�1s��S��/�68�%oS�+�,,f�_h�b���Ɂ��oR�e:!�D��U���'�I�oc�տr�5�g�z����i��$��VO͆�?�c��G~s4�YS	�@�x�ap�௰
`	zD��Ě���-�
��"n7�_Z��[6T��&
�3)�`�FlEYѵ
��/��3JJ�E#	��㆟��!�<�>��B6�pk�r�*����l�����Y�Qx=.b/�潳Br�p�h����Ϡ��\f�s���w�F\��L���D��;��ȝ3��&�k+��;�G�T�.*ˉ�3��,�(�����Z��u�6�ּM����q�����22�*�8��`5YS~�r�{���Q{���Q9�z�;�{��gK
��D�լ��;Za�-����/�Mf�旇3�E����1���6�%ü����������aE< �M��]�j�[�U�jE���.��{�6���bw�<�����L�#B�x�:!�&�W�F�%�)�̇���g�S� �����'��r�Q���U2d�J��q�~;O+Ut�2��a�p5�M����^�{���=��H9`�_���\��Ko�1�A����y�ť�e�ve�i^��y�f'��F&`�sEQ�TP#�쁤7�a��s{R�k�_��r��b�ӟ*�����p�;��ӽ�'ْ�ɍ2k�$mu#w^v:�(�O�|l[R��6 �D-)�tB9Xlb�#3��٪3��0;g�%�o�S�Fz	
��d>k�	t4|����o�E%A4�����=�.�`���+�vn��K����O}&���K��#Kp�>DB�� ���r��g$	��H�7�:��B��xkܴ��'1}<D��I�~	�^%��/��r�����Q>�s�I;�T��z��Ȟ&<8�H ����/�?�ݲ1����X��؆�r7-��\�xnl�g��O&�ʘ��3� hftԑDz���,y�6��J5Ë�h�H�{��٬t��?�qw�q��➼aBC��Hn/���Q�R��d�����,���V?��4��6�h�Ы��`ܿ�x���fм�I�_i�5��<�?Z������v��e��"������WO�N	 f� L9��D#WÔra��]@"ҙ�[�����陬�؀�Coc��v/)�j�������o�^�^p�p�	u2�#������D���<W�'�4?�zx�1����ocwC�V�%hU�V����J�f�g�ԩ�O���g6R���,Z*l�|<�I�EVR�	�ՀJ.Z,d*���o �_/���P�%LSQD���7 ����x���aL2�>�5x��5�}a�>D{׌?<���y��č��6�W� �ZR|!�"`/� �%����Htel����%��C�u(Ǯ�3�k�z�/1A�=*��/�*c�߽�\�6��H��P�*w�}�9'��9	��8'b\K-��Y�����p�ܭ4Gi�M�9^!M<�7��!��׵&:�g� %�u�H��1���
e�*O��L���d�s�s��qK�s�8�J�;�Jn�LO�7v]1\�^��EGf�1F(���&Bm�v�e.c�$בּ�]U�eCG6�}Ja��b���2�fF�ٗ<*8@D����R�i�a�qѰ)/�u/$�3��S�Ȯ��z~T��9`Kط�����Q���`�Y#�#�;2����7��`���2�i������o��=���o��D��҄sT��@�)ua�*@�~��z�>[g����/���>պ��m�Ƃ=�RcU�т�%� ��aS9������	�k����գ8��*=�L$�]��Z�h-
��$WgR�	_:�|���8��@7H�m���7C��l��z_�W�/��g3`��Wpz�T�����Z&�����>�,aޫ�<Kk���zC������*x���N@����`RDo)�{���{ ����LF� �eNkw�dA�t�6�g,�1��<��M�W�K0��JB��M�L�u�Uf��_jŵD�\�P����e�Z4۝�`3��s[/��5��c���!k��� RT������B(t�i�,z=9�z�����Y�)U:����'}U����H��(<N'�U%�4���8dc\������r�c�C.��Ë;l;�r��Gy�᳅��>�y`��
f�����@��&�W��:���́�t��ur�Co6��mE�rp�!�W� -I3��>�D_*F.s���u՗������AR����u-�"U{R�y����"U��&�B �~�e���[��J���obs�'֐�*˖u���"�޳V��� U�<�cEn��(���{ y�Km�ܭu�kT��Cʏ��;À���a��8+��@{z��c�]�9��� �;�r���d�R�����=�;�|YSzU�gbs;�>Q+3�bta�}��X���_���{0