��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��o�Y{NĖˬ���P/{��$�)f�Y㈎����� �9H$������,�-_6IX$�������ˬ�Zn��B�k��b�H)7b�WˠUe��Ǵ��A�VP0�0��{ߤ\z�ύᙉF˘y؍�����
����;����k�j��F����H��ja
�P��QK�悅��5�sʮ*q^���lF&��OG_�l�ic:ɽ�.9x��}=f��,aFz�:w�;��E��L����^q�j�k��5RBl���XN �\���a�Tr��kR�5�A��yQ�^f�n�ȇ�I)���;��~�xM!�ԧ=$�z�c����s~@�n߳1�����顭��*Ȃ�!����Ӑ�,��D��
z�@R���ڨ�0`|�Р�ڂZ��y���Տ���K�9� g��ėABĎw���"�� p�c��r9cqGdsA1R32���D�f	��Ț*��j��֔����w%s0?��O��!w1��ȴ���4��0�K����*wϒ��r��@|wH����@G�����}of�N�|�1j��!��q���O��oP�@���Z£v�u���?���<�󦏌�C���p�9C�N.���Y���?��&^��yg���emɵyC
Ծ�E��S3�[)���"��~ph7f�	�:b	s✾Կ{�a
$1��iH��5P�����e�����qyv�:�/�_Љ'�"��� �o恕+,)i���1�͋졯 -�Da����	�>�N��"񠩻�Q������c��ݭau�Z]�k5Y��!����}���~���N�]��׋��ba�;��� �5��6��EN�&�>�)��Qv=>?b9�V����sqTW�p�'g�Ӄ��3�A
��2��Y�2&
>�}���ś�4S�s�p,~�{�]ڟ��Q>w7E73�,M����9?��j���ː��-�p�e;�/�=�r/UQ3~\�Ő�7�դL����^V���7��gEO-d�]#&Bih��0TV�pܽB�u�r�p�>۾���K���Y��.U����p>÷��Q��K��\�^,6�I\g˶<x�2�z�v�\JAI���u�,~-p@���WR�=�Aeh�\����Nq�tF�Z�Xd�V���n1��1�y�����*���e�aX턲��4���(wZ��Q����"�"ݼ��L��YBf��`��`����ř�m��N�_�&;n����Lh�x$�Z]�b����ms9�*����d����@�R�N�����т;�u0��q����-�����A1�[�聐��B�O�����x���tt�Pؐm̍�l|5擩Ԇ����^�&�NҤ�mS#
5��y�2a���3ğ-.,�t-��.[��`�poKҪ�jLi�d�M�Т7�״_��8�0{+�f��1W�'2�л�S��2���n�O�?]e:��6��W&���WN8i���$	b��lKխ�����Un;�m�3��e^��>a��G�IO^f�Ȳ����J���e��U�p�m���3\h[�d�穵�)�[�M���`n�+ǵ�hs6��}�;��P��[�tՑ����"��@JNB��D���f�<y2���l�9��(��!�e�.S(�	� D�mÍ}�k��(^!3K�#��/�f�� X�4H��kr�8)�<C������O�����ط 󧶶R_s�k������+ ��V�?u�3	B'�Z`�`�M�_���.�r��Am2�<Xͱ���7�rq��D# M����^ D�g��Xd$0�e�q�����d��v#��$Ls7��`t��%O��3�P�l�ݒ�V�v��ЭG�%�BJ���
���zNt	e�������U��d�}$�	�,s�({��L(=�1�H���?��L͠Z�_wʶt��4�:������]ʥ�`%�H�� ��B6U	��L�ޫ�TE�/�鱢�+��$o�6g20��֬�|5��r]ؓ5��b�����s�.�W�J�-)�k���4HFDs$�O�CQ�릈�G =�����	�h���jX��x�X�E��%8�L>Rl��b7�C2x��K�NF?N/I��hs͝����/�wϨ��
*6#m�P�צ��ϋ��".�w�D�I�RJ���Ü��/���� ���T	���Oޕ���./},8�s�Y�~'��{����f����.Sr#Þ{4�rD?�6]�`o�4�����[��x�罖��JN�p�F���0W���E.͟�&*�G�f(|N�i��:ʼ^������t.I��\�d'�%=4�D�SΊ�io�Wܦ9U�h!#L7nI˓S�+ī�J1ۥq� �.��㬻�V�gL�ZNvL��(��l������#�I�i��� �Y�:���_N�'3U)Y^Ts
�J�	r��Ls���:6��[ǭ�r7��R%�U�ʘ�tf�����:��&/j@�L��uh|`,xI[b"���Rd��b���(��P���Փ��O�3eRV`/�.x,3C(&Q�t�z�+H����߭Ve�A�S��S6�+��H�1�Y��BiV�Ţ�<������XW���Qx2�!ؖڥ�e�[;D�s\�2�Z[�<Lf����M�ن�C��r��(\Ff�㼧e�~�N����s!��>������j�o�q�����#i���a��(z�?�
S�o��m��<D �� H�&�hd����u5��yշ(���U�9Ιh��N��vq~�Ɉ!��#jƴ��'-����D���p�
&���XD��s�o�A>���P�$M����ei�T�l]�;�n1�K^F�.o���ecI�/bR�b�������;Z+�\�M��w�m
!�W�)C#C��Ll}�)Ƣ�c����"tH��+�#2�QDm�<�/�<��X� �͚X���{��c�����:@I@�u<$q+c��Š����ڙ��s�_�<����v�oS\�l��i��ݵnj_,�ӗv�N䮷_��@���X_�
�
i�e��b�D��zS���jC�g:{^��1 d[�N'"�Yv��$�	�0������HSg�V�<��;�י��/�V�L
Y��?D�R!��7��)p��O+�\�z�I���ԅ�:�sY���EIA��7!�� i^ƍ�Xi[U���k	r/�G������ӝl6�v�����9��	aXE��0׿��c!p���N�J�V�R��(˒�,'�o���Ҵ4��J�G�vї�1n���	��Y��䟁��vgy�+I�сI�����N�����6�:N������?�W�(����5�&��R�}�E�8��`��e� �n�ZP�S�z�m�p��*��[]���*�R��.Z����+F̴%������i�g��^��b�X��[=!�ovL�PIR�w�˥�Zp��h^�HB`s�}
�a@�V�+L�H�#�w�����P����vˉL3���]����SN�p�5փ/���bj9ِTY�#v���-��`�Np�x�Z�ՠM����3(%$�<g������uROP6���}���@��{���I�'��n�Fn�]�$N��T:մ8<1>`�MM&�6>Y��;x�]?�)EQ,��0IZ�ܚf<~� q74%	Q �6���p�"�⹛/�oD�k��ȍEc���\��lO'��AN?<�6��A�2��<
x�6
��\�&U�=�AR�e�¡/t��~�����r-���Q}Kr�GqyՂ�S6���^�2�)�V�6Q��5�lm���Zp{f�>r�Y[�����Q�a�S�ژ��Ja{~.U����7/�q?NJh)��a#�[rf]H���R>���(�� o�2amy�M�޻Ϛ��5�5��P.8-����� ���·�LڵH�fV0��'�T�v/�"00����wDri�}y+�i_2�g��8��%���Phqs�a��pd�C��a"�!=��rS���|�z*P9V
��`1�1�.��>5Ֆ�\"�QǪQ��$P�+:���N��	
��*X
���*��
���<��G_��J��i�La9�}f��y���SV��=��3?��Wcb޵�C��� g-��V�)��g-3�VBY;d�.�;�@MB�:���j �K�t�z���!^���^s!��F'�R?��Iġ:���+Vy6�Jn�6��qj��U����@�S��)�M|������#+��
C9a�蛍mA,[l�u��&V�Ð�5Y>t�O@�L�	<���D���ڐ<����ƴ��Ml���*@�\�Q�ѱ'^�d�)�|����g��>��a�.��Z��L��/��_��&�[���Ԍҥ�^�)���.}ܥl�7!B�;H@����C�
����W!�k�[��o�|jO���޽Vt�|��+k�HǕw����k�5�ƣ�^���E�ۿ0������TK�x@�8��r��A���8�#p��=f�L��#�#NS��VɎ�K��`�?Qz�#PлUhhژi� ���H���ڧ�|����1S;2 �P5�H�
pU�$��jV�]���;�%�Qd&�-]��(��:�)#����QA��6ķ��D����L&D0+�p�C��S�O��x�
��	���,/lX"k��S�B}X�	��m�#���<���t�1��OBm�o��q��L�qj6�j�~��������H]��N���z�-F���vݩBϸ�e�p��{̈́޿�Jc0C�F��H� �V=�6��!x��>by��jTA�ſ�_��C滣5FU��:����3(�G�R��W�(�`2���	 �XՖE��|�)��m���A����r�<W_�xv�m̥��I����`�Vhup��O�vO����!*��h��zQe�-)�ȍ]�����2��mׯ�7�ym�'Ҁs��=�#��ϳ�J��w�@�v�Mp�/�q�߯���Σ��	�IX[�Ax�)� I\UQ�5��Ԡ-؄��"j��s���������X���<!�c!F	�>�^�!�@����1�$'�}i�ع�=_ H���JI�<;'@���$O?c��
��$|4�(�W�A0�VW{��p?1}�.�L,��]�I�	�P�Ê�����l�k<4�>諎s���ϜVXDΥ�����y��B2����!^=�2�p�0�S����/k8���H7�Û67͇dZ�x�_pw�b�@Hj�lb�rP��A�1��	X��m�����B��$UqQ�[�w�C7��ڨQ~���PO겂Ho�ya񡪣8�do� ��#�į�Em�}�f�:�p��n����
B���]�W�x=�ee��F�b�Y��Vܣ*Շ��-�9R,0a�^Z�;����R�}&�J��3�i̞�������uo��ƪ�@�/8���x ��>ˢ��H�A{h��_؅&NtXJI6�G'��4 ~�f�S��<�^h�s�D�%�$bm.���RD? ��P������]�l�l���p����k��L>��q/V����_;��F��Ȼ�1�`N���lڷ�#ۘ�NM@5J�x�W�)�E�*����ءR(�KB����@������$���� v��o +]b�?c��y'#^������G�_�M��Ȫ���A8��>6�5�����������(��	�/U(#���'�HݶG������Ktt���hx��v�47B���'�\b/��:��K����E:"X��o@�����I��p��fZ~�ԥ\�W����`�.�����?��I�3^�8�nk�^L�nl��Յu]�L�9�n��% �	�β��0�vy|yq�uG�]��Υ;�Jp��W�co<��:�\|�+��x0Q\����0�I a�Z��O�D�inK3kP��kH}Ү��2.�`/B��Ϋt]A:�Ϥ�q�8��5Jo�_���{�6�͊i���,���
t��t]�A���K"L����Jlv�"��n���w���� � ��}����A$!�/�}���aS����0y��R����{�^��.��	)ե�-�
vDV�w�Ia^|��6����n�| x ����	\�0��$��a�7�R�z}�D�lf3�-��Y�s$�&&Ɔӂ���tj2�ąQB�8%ωbai"�Q 'w������E���b���LF=z�i)**�oB}yk:�^�![��N�X�j���fs1�B����{G�K]+�AZ�1|��ޜ�'�y��O�a�J�����^T?���
����8:[Ε�*I̶�}@�c5����[�&1����_Л���!#T& �C=���Ic�$�4I�V�����@O)���t ������V�@#(��8��=�h��bۖ	���\M*2Y�t�9��N݋U���T䩫 �C�r/���Ӳ��J�Q����Pn_�X[�#)��+�|�Ka'wDO��A��ڬjwa�z�b����^|�+II.�H�e��y��u�g�#�~�6�����7Ǹ��\�Iu�m��� ���̅�̌9}+$V]`A�̞�_���:.�������=�7�P����`V�'��$�	��g��q��ג�t�#����>�k�i�fn�]R�-�e��f7CYE�X��7�������`�,lw�Y�d�yV�=��,��o:D���{q��EbD&!9�0����{x;��IvQ:�	�,|�_uS5oȨ�c�	ӊ�M�i�j�T�P�c��De��Cwa�T��_����5�bA�0���U3�7 �$B���4�U�97W��xG`��E�#��3�pzg��	k�Q�(�s[O	r��#�g_����ke��������J+T�ol�ڑ�ԇ�H 2�<k�>����~�>��kIx9�B�+�����8��g�@�a��.�2&bÅy��;�����/p����XT�4	�kY-�~XR�V��������*���E^�kS~!���K1��h+0�h�n�'?��rs�I��2��Q\���2C�����x�$P�\;���� x+��`��/�C�?���)���FDÿ�|\^С"^�W0bҒf@�IN,��C'�|^p�&�q<��O��X�j��{`(f.�t��+i������rfI٦߁S7���q
�&*�� [oV��ۗĖ:��V�?�A��Ā0��R+g��z0� ���9�3�<$C҄��I�G�ס8^_D��e|��Z��B���i;8ljŎ�a��xj�2��n����y&.���ĕ���MZ����%�������jC�i�G�����gc (�-��xjb�1�R&2���"#�,=�xe�Z�B�r#�kT�#rc�����3�B5��
�y��(�
N���6����/�Es�]����m5!l3��y���F;s	����yNb�_W��x�I����Z�����"`���:��̾�=��4o���/�͘��p��݅����e/��,��R����˲�(�*�F���<���D
�Ń~ƭWf��ݖ)J�Jp�w�"��ɨ|k��+|�9 �W�'�q�EjN����	�.�市>L_kuh��G%�<ڣ��-��]�ݐ<���:�m�Nμ�����Fe'��ܣ*�;���#|JWow!{������5F^�
Qt�{v/�mh	��qE��"G�*Ӽ��d���?��21A�� TԷ���Z\ώ�w�N��W�G}�;WTF� �_����8�x�F_'�w�k��_�4Y;?���X��g�w[��'��%ę�u��^ ���sl��Z��[� �?���J���ik�V��hՅ���#v;/���Dcm�=��"��7��!��6�N���"�@��wl�Gr���	�2vj}y���6L�G6𷉀�A��P�{�/��ya�9�95m<���c�?�ނ��Va7��7�`H���
&�����`bG���VH'�-�I��"v�&�	"̶���"O��P7$P�{�OߘX��W±��t�Q�ܭ�\�1�68�a��@\�sЕL�H��֏��qg��Mt�rZ6�L^��q���K�O��a�%��}C 
IA����Qo�UE����&��Ka�ÆjY�-$=�*,�YY�ThｳsΡ�G�l���D�/&�di�-�IE.��S�xr�K{�k��8�͐X��U.�o�����$�����}����@}�羟�m���I���?���ol�ig���V�	6�k&������R?���'ܫ�ȶu��,�Ƶ)�A��
����׿��vv�e�;�?���(���K/��H�yɇ��ѬY��z��EZ������&�&�iO����L�MM!��nIS��U{K{�-R�,�մ����ĭ�|�=�2L��Z��&�R�t�'1}|��������*�|EʱNOv�;�Ϋg�zZXxxٝN��7��g��*�4������֏=&���.��\��%���J ���R,O<���E5�jdH�$~��N,Hز@�K'Kg�p
0I#?"�<խb7p\�מݣ���[/6Ҧ%-8���K���]���v�d�3b��Π�/`:9zdj�R�t���~�[�$L4�]>�Ѝ�h��3<�o֓4Ux�-R�1��V]d�� '���H�cwNɎ��]�o�`������?�ʦ��Ln��x�L��wvQ,��isXD����,�����a�i�G[9gu��5D��>n����~���A�p �y.�R�H��� B����6��Am({�RRM#��rR�[��Dw�x��w����b�S{���;)������a���k4k��S�A��5�{�kXv�z{�$��H�'��.��3m��H�#r��@|��jv�SB��Fd�?���!�>|�^B�g�� �iNDz\���E�CY}����Py��]KK[|,#�����9�Xκ�<�U�����U+��yV5�l+pA�U#}�:*�џ�,$YJK�g8Y���?��v��}����O���:���򀟥�M�8�'Nv�BG��oF�V9i�ob�O���k�¹4۰j�+Gl �����,M�|_Y���q$���x�c���+9� ����]k2����Te��9��}����T"_�T�jG�PV�̍J~,��taD�U�8$W�Ĩk��F��wg��kl�/��GF�f�(R���l����39B�dg$&�#rv�E��ɷ@�j�����zd/
o�]��Dʣ�jZ��e������Nj�����*��s��t����vz:|p��Ү�Qل����P��,ɥ���	�u�#(9���%�c��Փ+���)Ê��	�Q��;�I�[M��/Ǜ�|�h�L �d0�_�[���4���cQD`���C�<[,	��0�
���|�^����V����,�?��<��В�`,I����_ �o?Y����OE5��+n��δ� vk݋���m�1�M9�R�J��󤍂��,�*��0��Rm���6�9��qA8��;��%����J�h���2��޶g�M�vIp4XTvAl����_XB�Ș�r9�	By+mݷ�V�t�]�C���
A�I����]�|L��t5��i���14��8!B��"a�NSN�@��&���u5j��HȬ�:K��49|�kA��J��ғ� A����@��7w��/�������(��#)�0D�\�4�����4��`n����i��59�k����[���QpF���Nc�c5S�6;�@p�KQw�.̆	���D��+9�8?�Z���£gM�+�.�]���H��h����%���-^���T�~��gW�͋�d�g"l/O�	�Ƭ7:[勱��t��'�|�: ��&��k�L^>��7W8��rS S�.Il��8���2VXGΡ���FB�F��=�eF����2D�����e�	j��^9�t�f'�W��n/߇��@̏�d�˛]ǐR�x�r��r�#C�~Aô�[p��$����лV��{!U���b�>N�OD����>�����LXX�;_�(&Sާ��FJW�^���ʛ���s>5�o@��Ԫ�EPXG�6����t�hj���#����Pq9}i@����[PQ�T���׃�D�W��� k�7x9ckL[����`s���f����}�$t/��ɊItӕAX5������͗�٧��s��*�+�Q<�x������e�	�6)Haep��P^c�W�����03�vA�;�b��vG7�����R�Rn�	ٝ^k�ř�<M��w��tb����Wp��-
� ���ަc;�A����K��g{��3��섲�;�l�`�@��i�4�9�@\.��Ǵ? A��f�?l�*��y�j�p�ό�P1't����P�;���[�m����+*�����������Ups5h ��K�[T;�F���}a����ڍOO���Ń�P~�B�'dll�3J��/h�f����9Af]�]�-�83�O�z0͛Ǣ��q��Q��o3�lxVOY�l��7��tA|����;ƿ�Ϩ<�����r�W~��❪F�'�/���K����,
멹����k��{#=��ʎ��!�"A�w���2"�ݢn�싫�v�gO~���e8|y;s!n��+�>Y�ϥ�i�y��	Y�j��n��f��)�XH<�F����ׂ͡��9t�a�t���	�ߤe|��;v&~��8:S�VS�<ҕ(��܃N^�3�eW��t�\6�v��+��F
r�_����^�M�E����!W��1�Y���r��ŧ4̽�6�QM
�0�n�q��p��e���SjI�W� �A��f�y�����?� ճ�����ǕF��㼨�]��a��Ze�8)�'�6�֩t���R����=��ǡV��鲡h�')9�-u�n5����$���""#�o�2����n�^(��dDm�*ȦV
�C��t~l!1���]�^�ʒX)�폇���/��p��P���2#��vVK{�0�֜KKRBA�����Z�#^n��̻�g/im�h�H%�('I:�p���i9r�H��r��}P��r��z��c����_�q��͉�j��C�SD'i�6�\{�H��+dB7�7�� x������oI�q�rKW-
=�w �C�jo�}�M��47\�RU��9n�����@O��H���΅ǡ���,U��^>��,rd�z0��[��838�T�C�Ё��K�����yi�S$�Aܦ���d^\4پ��O�u�3�r����N�h,Ĉ����Nsо�y�p��~�`���G�ŭ�2������i��;j)����p��G�&E��#D��+Jw"�:�03�1�����^]O"U�t�؃V'	�'*g�:����ƍ���M�z_�K�����HZ�_������A��!2 ���w����L� ˲�;��n���WVYt�v��״�hp 6,�!�m��B��66f��U���m�Iy9bN�XF��� �)ߏ�8��R���ge����Q��ދ�n*�c��f����yJ!CUz��e�h�r�U� �ȶNC�@G�n ���g���V�d_8�'cjԅ���6 ӳ��{��W�]�S���ynj��u���0���.�S�W��� �UMz�@?g%�]L�����!��(����3E}���6a���F�MR�]#���_��t�BW�W���]�+��@��8�����	�e��}���I*��Ǹ�xԬ�1�3���S���|�MV�e������f���"]�����E�a�8x�v��
[^���YB�H��p�N�2V�F�Pv�4��z#�����Z��!�wZ��Gi������-@rr�V�sC�f���B�|k-6#B<m� �׼�gg�H�Ә�Khj�����C	��ۓS��� ��gj�?�(��4$��$P�,��M���ɩ�N�������νfzx�\H�wGMU :�'9��� -��K���i�+���=��`���Ԣ��Ì��W���葘Ŀ�oXqF>�֠TT�i+�p�\�,;/-h�:7d!���C���4�x��2��v����,��[#$f!�[a9s���M���.�R5D#UD�gT#�x�>���jG�d���ϡJ�ڗ������鲯8h�9�(�琐������lGxs}�eT5�V3���
�0K�s� ��~MwV��b|l�eJA��XO���tZ/!53QR�f���q�Ta��ܗE	�C��%VQ�(�5���
#p�?��wa6li4��A<���Ɓ��-�/���oF�Ҳ""Am?��� �[��T43=eק8�VѴ85H
�<��5�D�b�yI�=>��c݁y-!}��\���W�>�Ѕ6�F	M
h<��i����yH`>9��:1e�!?K.�M�p�׃�[A�[��N�<�D�e6���gdڠ�"	��0CP]`��]������[Z1���i����+��A�/����4�C�[�YA&�"^ܓ�L. �y���xN�z�/�,�X[H�H���-�ފ!s�Sb,33Y��L�������-�."/��k
�t]�����T"A��DO�{�?�!y�|_��>jid٬�����CRi�W5C�"D�kFW��l�3+M�	�8w�_��;���,�$BZa1ݝ���Ɲ�6��'H�# ��*�v32�W����1�#������LdZ]$�MW|�������(>��'�o�md8E�F]F��R�P���ra�]q��P1s0M�۽��3J�^���=�s'Y+���3��i8�wfGR]������pUZ��wU��*���N��E��_��8�C 7�wI��r1�I=���a:�������І�� ���{�:�~�O���h�o�Ky�$NO��t��[�Z�[��~0��-�[��4��LM��/�X%z��y@}�A�rt�8���m[+�yW�S��'Λ�x
��
���1@Z���E>���W���&�67JX��~E�S�� !�B��qfGh�E��s�t��_cCmy� �����jMNQ��1��UI���ײI����QQ��Y�����-۟O�j�_�('������">vOx@��a���6�=�u���~q�eN���ά�9�)6�]6y����9/��IG��na�rv3�d{���mb��/�k4��W��ў�tz��yz;�ho �>��YIΙ�c��l�뿙 ��P��D�՞���:Q
��������]��x��O��!RM��/MW_�-�L�!rp�@ǎ��2��?C�E��!�L��7cn��O\^����i��|}&�PP�~O#�Pʠ�'�hL�Iȥ�dޭ�����G��bB;?G���U2h�jY���oC&��,)�c�,�Ki{�F�Ѿ �ͧ��=s�=Il��`����'��"S���.��m�n�ǒvl2 ���Ap�l[R���
0.�:3B��k���U����+��r�*-�����"j���gH��b���#}��uJ�R�K��f#��{�u9R��Ɵ�
y!*�0�� ��?���C)h7�L�4A��^��sO6�]	��^o���a}D:��
?] ������H�t\�$w����KnΥ �;��dg+=���.'���[�����>r�O۟zA�6�}�J�+�. w[\ �Џ&"���^�(j�h��H;���F�o�h�uO@��b؁[u�?(
�r<����C���̤�3�,+2Q�Ǐ!Ўr����7�C3���!��Ϋbpjz@�3��^����5�e��C��a�#J���|-�R�"e8�'�_C�ڸ.QS���RW�tr�H�� =K��Gk��XdB�`�X���/����lc1B��	��??4�y��l��H�Aa4s��H��ms�ٝ����c	�֐
���+������E�^���e{� ��p�Õ%k��Pۓ�Z�LCD}?�s��t�y�
?������&s%�E�]�d`����,ڦ(I8�x�˓B�\��e���j�+E7{Z�$y��#��E2'�s�ƣbF����؉vN#�m��Ww�ަּEo)��H�U�?�b��]2�y���^�B�����} �,�����S�q:2�ɡ�����Au<���R��<�0�|{�6��*��/v]0��%gr�F�'/ ����]W�~yzCv�ώ ��ozI$��M)��x���Iʺ�"(�������5�nzb���g ��]��-�[߉F`LȔD_*\TSME�1O乣�К����7��߫�gT��P�B-��}x����ÎڀV�jS�M#�  �w	\u�AF���>y˜����I]��gӋՆ�����MfkqN
�,햍),!�p#G��	=d5�_��'o|�"މ*i t-�6wN/��G�1R��2kOw��g�7Ǒ�&���4��9lqe)f�ǹWBo\�hh��P	�~�����X�H&�rpW:�̞�]���2	aW�i���{��������C�5��i}K!l4�7�`θ
0����0�`kq e�#�1��eu���Sa�a�\����\������Dn�E��Ӕ�j�P�bsZϔS(U��%�y4o�>�<X�����X���f~�g`��q-g%�q�sY�,ҽd6�yEy�M"�,��yu ��j��>ad�KI<Ϫw����}�&�/΂����^2��w��d�"n���}�����κhm�Im�8T�x�x�!�0X�u��]\�=t��~JuD��7E�x���v+��c��y����u�I's �W����;�)N�,���8El�熄`uk��L\��RrR�>��kzE�l/����01�/ Ld��$Ib��`\�H�en�ښC�I�e�hH�O]{R 
20�7(�4�YK29z���y�j�Lҙ��&�����[���2l�䆞�s�
�{���� ;��z����ϟXG۸¶v����O%���k�2��d$f�ߍ�����c�z1�S�'���b{� Q#������8��n��5�u�9�;���N��`F�l��k�)�(�D�c�5����Pt��n\�ۇ>����?4�7�\�Z����N�.$R������x�#C_BOxC%1��^L�3]��K�k'��?y�Q˃�j��`��~I���eT��ɖH�������7(	Q����Za4֚��!��1Ό�|�I�H��r> �n삍N9���+�8KZ���Õ��)`$uup��_(/8`������U���3b6�^|%O��H��^�iwZ��s�R�D3U�5k1�^�^oZe�ǅ�%&���c��+.�C]ܭ���uk����櫕m3�i�?� $�!�}��n��0�����,�ͺ|E�J�Sd��"��$�D�҄[�mOs��}�/��-r�~*���$(������=Q�X�O:/2K���r�RZ|�S��=�^�S^=N�Y��NvE��Q�%X1���}F��ź�z���)
l�<ZG�Nx��\� `e����{6�&���#(�VIyg�s�2G�1��B��?�Qht4$�Ks��>�[p�D;q��2�o�$���M�_m@�!�,���NǤ'iRI��3([� `vѨ�YlBf�t�x�72�����$�&,Y�y͏9�1��5`,0V��ց�R�s�y��#w��W����B�>*|�s,� I������3��l���&�,��UE�ϼY1Q}��� E9U���a
3Lڎ�v\T1��SM^j�rEl+� Re֎فZ-\��T�� /0�6�u�$3��`�0‪�X�c�ChL:�	�rK�B����aO3 ��dc�����$��|t.;��teUwu����1it���,�Z�����,�b���L$�/~��z��y9)�N��-�|��"��dSY ����w�9/&q��@B��GQH��LV
���=�R�=z�D���+�aF5J��*M��/ac���PH�'�Ρ?_��4��4kG�j��{�g����E0�0#��>�<��ts2@��0n(d�<l��1+WZ�_	u�=��~�g%�oɂ^���0�CY^V�ڑ�=�~�7���+Î������s�?s�Ar��No�^�Į�hŝ{���ӈ��`�";f/�2��`������Y��S�����]��^��i��9k[Sxi�\d2���DAū#u� P��GՓwnX7�-���5SZc[�8}M�^��� Lj��be�"�q�t�:�?�0U��� W�����׮�)q�̟XY�V֡j?��<Xs^����7M��
�n�jh���M��JG}�X�]�d���?Ϙn������q�z�B~(�E|�V8 �*-��4�� �L���(����o1؛��QA=��`"i�A��Z�O��N5z��__rY�#�t��D�^i��D b�>�?i0H��h�ٲ�mR��/�B�<T��22/Oq�ܼqO�	a�]+�nbgdϺ��"���M.�D��A=X�W{	`?Cs�L����]����6�L�:0�Q[��z��f<���T���/qK)�`�)m�}�6dV��'�+��C�ר��F��<B�}���H�M.��[B�F5�3���	B�y���ˢ|�thVk��_O3r��MlhuU8U5q��s�96�qe3Ar#�g�3cOo03F�C	W�&?5�������e5�-x-�.O�<�l�-�V�u��y2���exȲy�:т���ݪ��E�|냢�� 5��}��7��Ł������³�>d���(n0\�Ρ��n�u���<��g[�h@V�#ݥ��P����(����Qek�%�~�Mf�U:rٚ�O��3�P��$�&��2��|ؼP9�{Z��Ygm� ���E����ӛ�B2��� T`�
e\�Ђ�B�����4%NR������m|Hgem
�)�"Z]��s�C��+ql���Z<B��u���"��C�f��'(��,ï��0t�1� �\�g=8�CQ�3�A/��</p62=���X�)Z�6y2�S� �V�����Lk�!�n�M̝b�l;eV����s�i�� ���M0ix8gA��ΖJ/��h����TW��v�,�İ��_8�z��D+�y�d��J�I��P]|zq��.c�o���a�<���\��}����)�&}�͠~أ�v�ӵ�K��x���,���C쑫���(�{���[b�$�1�N���d/����U%���raC�6wʌ�s��6���:���:��;Sro���J�?G�i��_(u#8��`sҎU�Z *ny;@Y�n=��꟦���~緍cTL��r���!kM��{���i���i�\6��婯�G"�Q�)��@,a ��b�۾pFU��@���Z�(����x�'= ��B��hK�
Q/�V]��w�D���~���a�f#����L��i��[�$.�>P<{FB=,��Ҙ�n�ۓx�CN��kc�h��r�؆R��1����ׯ�)��ɑ��dBx�V�	���=J��ˆ4�5Ax�[�*SL�������%��~����[Xި�m����qߤ蟓
l4�L5c/ճ��Ͽ=�wZ��@˕o�M��K<"-�@hz�xۏ��Q]t�����Ρ4����3lS-�b�7.��ē�t6��O�CM��5,C~{�P���
��P��h'S˜~{M��v{1��-�/��b�Fm>c�����2�3s�7�S��i��FSMɐ�b�7C�����`l����W��"���Hy���7�Z��h�ʯ��YfG�z4yH�}���J�9�0�d3�DҲ-����!3?#r�x`T��x�/'�[�ǁgH?�M�w�6z��T+q��+!��EH����]���q29�\���	���rE���7�9�J vŭ�rCj�
D�N�ڽ\���M�,}y�9����x'�s�}�Ӯ!�v�FƪlJ�V�T�~��":ݾkCE����}��kTS�/����@m���eg����5����}G�3W����oH��+_���"7�