��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��ov���CӇ%�â��Iږ�mG"��?F������J+�އ����}fk���������C6V'ͷ�m�gG��"k�� �K�!|X��>	k�n�$14�Pq@�d��o}���VV��b�M[<rU����'\�7:{�Ws>/Z���O�ʹ�k��\~sH7���G��~�"����]P�F�G~f�c ��b�����z�y���9��`�����U�c���OMh�������o��J������l�NY&Y�~�+S�>�~�����1��}�: <`��gk�#v9"�o�C��&bb�D/�^v���L�p�G��%���tj��9�LF�~�e�s�z�_���#)
�R	�'��^����]�uꃈ�n�J�#��r�D,Nl�㤪?#�����\���E^j��M�8��h�%D�Vv* �g��J���l���G����{L�Tv�A\�4d#x�~��w
���!���+�0�8�p-q�nŰH��1���1>4�Z���6͜d�=�iM��b�g�s�զ*���lsk�ұ�f�l�C��ÝLJ��<���Ư郔�׎l�"`�[����kj$--r��@�l��u;fp��e:��v
FM\C����R�����U~��@���*�zI�������1��{���f�Z�C�G
�U���,��o������z���C"ý��������z�Z��zji����XOJ]���(�x-�o���",d΄4��*��Z��|&Qķ����(=�P��a����}��A����z�������ww(� �n>{�kU�`,?��n�J�gք/2х���X�`�wRޮ�F=luE��u!���D�f�"f�O]TPx��M̌�<��Qm��z����N�>^	R<ǯ�Ӻ�qHFQ�l���6��D@i
pִ�mȣ�F���5Z�2�� �X�S.���w���ȼ.��}!?&�����s��F��w.���!�b5b�MB
Z���t��t:�4%��>���ّd)�I׺�0¥v�8�ai�e�7\�8�cA{-�U?{!mx�O�,�״�zk��K}��_.�S�	�����7�#�f��8o7u�	 ��
�1D���`��	]c��@�n������Th]7��O���L�e��\��Tﳯ?����CΤ��wSE��Ņ�s`Fڮ�٩A��?�KB ri��[!H`"f���e,9.
��Z�_��e��dz�Hb@?��vt"f�!�.+��s�>�R!x?1�=�D�����M4���xDL�/����Ly�{%(�6pOvzE�+	��ǫ���|-+��ͣ>���&GS����xE#�\Nl�q���č P��3	~����S� g
���r����z�9{[%�4hR-Vj�_k1�zN��	���i�b�y'���RoS��(�H��:��kt`�t�߽F!�={�*�|tӰ��\���ѭ<zBlG�����W;��:�q!�-��$`I,u��v�UT.^G�:��(U��G��]��-]*`��s�>�t���0zMb(Ɓ�@
�4E��c3o�{(=@|+)[��#Ey϶*�R2�uGMo"J�Ѳ��%[ Fm�l�Aȉ���]>�R��oF� -4;0f��eI3���[O��b�5N;��!�������[���ۂQ�7�f��y7.e�ƿ���p�g������	�qC���̡>f�5�7�5S~��E)/E��^�w"�F��4f�׼#W4jA�#�F�p�_�+��� �Ļ.	�W�a!cO���^~}�f�cX[],�)��"�O�؆4��z>� �	8�����v�v6P'����I�v���*��)��1�K����\i7��w���KT�l����)w����4�v|R��?F2SPkO��]��~S�;��V�
nZ3�@�7��Q/���$ӭ�S-���'�o�С]]������[)�;Y�S0�U.Ů�_��5�ә�����f�[D�X������D�s�9�Qm�8����RP��y������n�u�����^9K���S�W�n�I�F%�bx��.���l�,z~NuQQM E����x[͘Z�l���{>��8�������9O��T�!�v�g��f#�uX1� p��`����H����e'?s��4U=��/h� �;�+�L����Td�0P��m`��RK"0�E\�QJeDd[2��Gy���|��O�]_��)��l��˛���cg�{��&[4�Q�`#�6���B,Ot����XG�樶;�;n_js��p���1O#ճT��Ʃ��$Rܪx���H���l�.��,�����v����W�.����0j^^��31Ņ���b]���T�͒���6}�(���|�#-%�����|Jbp`�!�M������gwJ��|���F�ԛ�J/
��">���Ws�x�>��7�F�?�
��{�)(��AcBQ�6d�6�C�F�����c<DU<�����hP~��
Xa��6���9L<kE��Ǎ�M�kh�@�{��e��mVu>�����=e:eY����Z�ĜD�}�fm���.ưa�,`5r�sԃL�[E#�
�I�,�V�a�`�m�׼+�{��/�-���(�¤nYШ�ͰѲ�fZ'�\�nwd��s.?r����W��@=$�8��-��޴��\ ���=j\�k���V�9�)C%�2d��Ԛq����H�E�+!ؤ`�Sv��u�q;48 ^b���o6���.c��1�ј�c�`=�~}i�uRrȂUD'�����]��.cĐ,���8uF�ςH0n��û�1�窆��VQ���E��OTv=�f���i����f6��$�/�j�5i�� e���~k/�]��@���v�G�ë�Q�a."+�WL\s��_��8:�0�c��� ��"���F�9^��B�Ҧ��H���n�R���#�˵6�e��sȇb�ھV�]�94i<b�'O&it�����jʱk ��'I��� ����}%�B�\f/����դ
������s�7�����+�������[��R*���_.(?�u�U�����Xp`>�U��(.���mZ��xޙuj��MGQ�@q�k��d̰���.����EM��Hw�x�ߴ�"$͑Pu�(�y��3��
�<[�vt��]����,��g�7o w�&}�du�Q:�9t��yҪ��}���9abf��C��p����;��B��$����i�r�7��^wh��⋻�Kg����eL	t���������R&�k�h#[�Ė�!)V~��2��R���Wt��,���L���4k�=F�Ȅ`��ɮfՎ�
���w��H^*+�<BkK�,�?W�Y���K찾0�ƨti�E0(�snVȬ��.�� ?i�}yO9��2��61��y^����5#f�5�m���	��y�M�:g��2�$��oX�`X���ua��r�&�e����(mj@;��OL�3��I�4&�Cr�7vu7���'�7�#�> ���Е�����ѱ�h�e�3pП�����Mi��H��>&��("G9_΍Q_d��_�:��U���T@QOd��X���#��N~��FM����8�
w�����L��>�s��!}�}�ѵ,6�3L�k�G�s��>�`�Z����\�5S1����=i�ǌ�9cA���d��T�V��E���4��Z���벿�hX��ݨ�>�o7;��Ӂ����sI��k]pH�kf�b�����V2T��sg�="�������sS}	�vE�K�f�G�%�7KEǁQu�����Նs�6��eOv�t]�@��7^u�Ї�dP�	�j��,�q�h��\<K�|�,\���_,���Ik��	�d�k�W�P=�V2+�D|:3�l�Q>��8���!ӯ����>��O�w!�g(���O��I�+�ǈ6�by2E7�f���]�x9����^��,�p��SfnF [�.���+���" z���ϟ�T~�~]<ڣ���X	�1) �ju���
2�p��o��K9Q믢���c�/r���p����o�z�)���N:�5(8(q�fԝ�=_3�T�N�T��|��p�Y���ϔ��T}R�0qy�jM:W�Zu\YCZ���箨���m�(��X?��ߜ_�ŋ����$w�a�WNcg)
p��S	�x�k[Za�|� JZ�8-�V8�j�jd�*	A�����������z;YB �S~�x��CrD ��|��ɉRM{ 갮^ �wn[)��_O�J�Z��U���z�p�ꢽ����A�2V��ؾ�d��O��>�����j��'VG��߇�=J,c97��HOmT�v����&��?[z��t"nW�U��r�Swliq)��8��y�!��A0lG��b��S����H�����	�qJ�Al�U���7�����{G��`�i�a=ti�����J~��7YY��R�cR�P����OZ�Tמ�F������_����]�p��||�����b6 :U���6<[ʙ��]�_Ъ!��h�*�|dK0��7̄~ }��8 1
2�1���gwFkt/c5�dNn�lE�Gl�jf�8�0,\���u@p"
Ce��*}�n3�4}�QSۊ<�;�s��͌��#��b��v��L�`��0�贪4��V	8��V��{1��������g���ȌH.��7�I~򌓱e&���/w�U��T��q��3���>i(�I>_���\�\5���h�qvJXuݩ���:`��<G�����R���A�K�����嘯P�kw�jz����{�-�:/l���+Ԗ�k�`��0	�ȭIo�zЈ�'��T��I�)��+�I��ʰߒ�
��?�k`VدJ���u��]�+�&�c�&W��t� &���v�z��U��ɿ�>�|`�)І�w�#>(1K���u/��s�ud�1/ �7�SZ�6᧻�Wk��ԯ-R1�"IQ;����m�wʑ-��$=أ��J�8�r˲r�I�	�L4d��Sf�d��W���� Mg�x2�ۙq�np'p�^�O�Af%H�����`jp�Q*gn �+U�)��H���k��F�#z�rC����0R�$f��o��Vq��q�SX��M[b����� � d�$Ԝ����£��ag��/�uiHjDd�X��w�đֲ�jb�O3/��#R$IբF�I�,% Ś�3����eC~4e{B�M'��H��m��n,6s�"�];Q0w��u��H}��}3@�Ae�!�XxV~�ϿMp�1����+�5Ʃ�YQxˊد�}���ܶ�����?��uC��ܜ�.��z�V���])���A~�f���e98���yn�C8�@S�B�F��ܸ?����MD��_����NTjS[T)���D81�0�2��b̔�x)�T�o���!{���V�uҕ��}��.}��n� ���ܰK�;�A���V��oD�������c�����F��|JD��m��:��=�<X1�#)\����;Ï�� _ޱ7jT(Ԗ�'o��)[M=d���zZGRqQ��M�Sr��2S��Y��W֜F�|�u@��U�]�2�6Hh�Xr��N(X��Z8�h	� ��2iq<�n@2�Zr�q�G��:1�?{b�C���RJ@�h.����z �T��
1d�h�F3����
��}����؆G���_~]�e+KU���L��fFI����5g�J���>eSn���*���PS)�t�EI_5}6�{t� �<67�wM�M��EJM~)�pЙ�_����4��+:4(2��hu6��Z�L�ǋWI?�NB�jW��N��}5ՎF#��� �WqU{�C8�ʀ�*��q=���Ѧ��_��=
g;�H���I;	o���p9��o�x�n*�*�.^�cq�z�	:���֧C�����ms���y�gOY����� �*�7��f��	bNm����Z���ͺ�7�+���h¾	 ���b_�Gu�_,o�-���@bw���s��L���2fc��$��NKd��/���D�3�� ߇(���<@�$;,D
f�&^��|t� �J����a8�*��n �2hk�l�n�ӊ�U){���.=R��Pj�G��� �lx5qfr�^A\��F-�=��4��Zw�t�°Զ~|�(���j䱻�z�LkC8�w����5
b���4��±F�j�/auj��ޏ�R���B4�ö�pp�xiB�I-rO��{���(����]u����ĴG����9���HKm�ʄ��(��E�g,U�[�1	��)d�
�Q3aRQ�p�
8�rUw y�����Y�t̋DŠn$p����ZA����;u� ��*Ԩ�*���ϸ��q1ӏ+������F�Ҡtk�n�9�{E*\��h�?�����L#�^�������I棖�ݓ��9`�(KܻT������ο���*����;����T�N�"f|c��*S�pT50���]��!�PJu}�0/5Ζ�hF@��Ws�I!����U���n��%��X�����t�$�S����Z���q�JT�$�8}/�y9z�6V��U5BY�㉝S��~��lq����L�l�<3]��Mf6�j���*�ݖ�+��;��W��`6�M����n�|eX���>���M���
�K��W8n�}Ё���X��Y�~�"��]"�;�٤����5N4ö+�C�?7��B�������[��+�o�����A�"A�{��*�n�8��� b���vE��PyM>�oa���S{$u�|#�J1�7lm�1oݲ��4�@����aҳ�C��	�q�G��f�s=*��~@?=�A*�E�|a��'�( 3_n��~��JJ]�6��L�k��Iψ�eJEwJ��QA���*��tO���w
�����YC�tR`:�J^Ä�,^X/mR�٠��^�4%!Ψ�"��e`}�C"#��3��m��쪨Չ���ɂ+�?o+�R*���&e=w��IF���'VV���H�"E���O���"����[6��C�I:s_Cr�/����[�"��ZS7�i�(֔5J�C_S�Ț<G���Tu��8;��W���s�p!�(g�8��n;YWG���ђɬZע��´d�_�c~����S����XMd��
�c���b/>�K��x�Ѫf1�}Ɉ�pV�W��C�@ �1�"��		��2�����l�7��+c�pmu4>�	�s�%f�.�Y&�`��`����Q�F��/��z�Q����s��ZA�I��=��o��ң[ޏE���.F�R����x����I�ċ��e������9��/���˲�mW�6t7y+�Y����,A>4n���s�_�������':��v����th�~�'%�^�\�O��$"�}[DkOwt �ҝ'S��2f=�}���P�����~k�Ų��(ׇ�B���<{��ll�_̓`=��%i\dǂu��
C3B�Dgu(ӧ�f��$A���xa.|�Q9�I뺈���갮{�EI$��x',;�G��r��"�Ͷ4~R�pN�>��O-<���Y����n��N�	z����ݐf[��g�@�:��od��q�Np���p��ݚ�A�+gI��A�v<[�W�S�$~�5lyێ���@-����b�j:M~�K��yp!� �:Uu�
�鄠�v�Te{vw
'�4ռ��H|+��2�%�^�&��.�n�M�{ԗ6�m�t6���Q�=���J^�HP}�*F�:��{�[<#��$}�³r	�p恻g=Q�f�లa�_p�͕cH�	n�1�'�E��N�6�E��̶��w���R��Va'C���Z?��1qUzm��%���U��ҾĐ�h6dI������΂H��ui�J�l������y��ÿY=׶��q�B	�,�Em>�2q��p���ބJe
�����!aɒ��i�����j�S�E��+���{�W/Y�tH"�l?��Ŕ:�kGk�Ō�>��0J[���Ò_{��	�^3�����"����\�{�l6�'F{Z��<}U��%��gKƇC��BZGNw1&��]��o�⑺w���Ք�����0�z�DZ�lK,Ҫ���Qſ���ɹ���=;�z}m�8M%NOQ�J@|l����lQ��4r+U�B��'%1G���/���UD�`��t�=ee�QρDc�xzqB��uHXr����j���	����\eΤ7����֠n����p	5���~��.�Z��=nbk���?Nb8����j��Y�;��F:�v;��3Q3a�ӱ�GltA��p�t�v��b9FQݕ�X�ܶ�3�j�������*:��(���~M�Z�D)GxI�!0������	�ٷ�#ҼI�=�����a:�0]Ǥ���뾱C�<���uz���X�ܖ9'�яŪ���xױ�n�/��|�S~�K�T+�]��^�n��-�3���(~7�������o��%0�ؽ�ӹ�VO�2H�/]qg4
��ݑK���f�e�GR��z�ɋ����~f>��i��N�����K;�_��G��Dy�f��-ݴ�amp�!�2�	�X�˝�60����ή�E-WA}�V��D��b�u���h�;�k"�M��6� �<rL9/S�s+_0gO5�J�DWB]�Ir##����.j���k\�3ȢA��$��fc�{�^���������0�
�[#L�x���2K�j�YɥX,W��Ŀ�3�W������)��0�~�;F����'If�\v,��@�k{OŞ�ӐT���4,Y��I����1�˘-��,5��/�z�}b~^���O��O.%W(E���G�R��}؞0�9xn������e!U�[��~�X9rhQZ����<,�eZ�ỿY@�!4J�ѣ5��7*��ԝ8T�����0C 4�huTX��?Bt:1D�ߪ�?�����I�8ҭpt��x׎���"0nn��t�<�'��0sW�p'���%�Y:S!�w���B�^W�|�a�(�k����|!��P���󉍊�ߦ{�����,���؅��j^���<��>qҏ^~�� =X���Bp��e����t)���(�u�2�ݍ����鈸����J��A�)V%X����?�}9�,���_ٕɒ��ɺ��BS��?@~5���~�P�v���HR��u� �Fh]��p���<+�J���A�0��7����I��lg=5'�O��ڤ�~f�w,���W�SW/J���i�7"�\��óԌ�l�4	���F�;�����O7T���}�[Np��D�2���`&[��\�2 �/%�L�}1.��b.��S=x�SɰMBx �c�����1�傐n���C�ߴ�j8D>-�i�I �Hz�~?/�O���/k���!��Y���G`hk�;�I^p�t8=`r��'�A���Q[��Ѯ�?n���%�-�Ó ����P����K~N�z V��k�5���Y*j9Si���\Yo^��AUى;|�?Ղ��9���ߐ5���_�,�;KF�c*������J8�C/�"y`
K�v[n���l"��#;����D#g�ԧs��g̣�E@��)�]Fb�  ��[-(ϋX���Bl�A��őY4���@8���XG��Ik�ݷ�w)�e%�����@�jfZ����tK]'.�>U8�k>��KgN5�J�.��0�oʰ�
t8�����|��G����%�!F�,������zŌ�H_l?�Q�e��j��)N!f�2���7λ�%��a���'��2�R�FO��;��_�� 
a���l��M4�v�W�2q�zI� ���Z(zH������ico����$���)�z���Ǭ��=Đ�w�&�*[�w=3y*�֟wa��i�m�<�k��"�n[��.��HG�!�2�~�P���mhf�
��qo�.�A�r�&
�/��q:*�k�Lz��h�ly@n����,������ٿI$'�@O"pYa�ة	�^�0�)䈶�_�$���/�E�d��U�����W���H�K���>P�.:��0���1q琡bP��8��f�}y'@-�Cye�Fi�F��@��&D���(��T�u��o��������cz��I	΢'Ss�}+C~t�=��sv�U����y�>�{ך-&8�c&
������_氄��&���W��B�5LYZ�@Gb�4�J8~F!���X�S=Z��@i�5�b��ͪ��L^�6��}h��d���H��`8���3w��E�Ֆ���-�p�Sҹ����wu�B�fFU�:��6���yc����ͳ+'����='#&�����dWQ]'����V���-r_���fNt�O9�3�NdQ����Һ��S����ҎX�L^=f	��I���*��%ԓ�l�;^�Np߫=��ӭl#(�ďS̐8����p�]�}�N'%�����d�=A�n����