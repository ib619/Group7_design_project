��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��o����\�����:=��0XɽC��1�o�~��V�44'����x�/�s�ع�ݤN�6mt����M��d����.	��r��C{��0l�d*9�{�!ߑ8�p�q��}nj=%X-�_�?�����q�w�?<J���t�>!6��������q�Y��Ⲵ����~�<��t|�:��	��	N���:lw��tf���#-���X%�w�S������8���-޴���M���sȭ)�otMp2��A%Q�$�yR�)�� *�*�
�L�ޥ�d[ַ����1����iVb+�f��Z/��n�%i�c	V`����T�q6I�Gj5�C�]M+�0�j�!<ZP���2�>��iZML���i����f,���ۉ\��f�L�����S���B�Y�yf� �(���������(K^��{�]J�&��	��X���A�wl��ߗ�dꚆi
i0�9f���~�(5^_�7���T��݃+'��Ym�<�{ݗ�tS��[���)���w����&gH`G5��V��l���SZМ���"����/�T7DF��x�w���MvEI�r�1���q�&İ��1p+��6�Ȓ���E���'t��Y�K�PK��m��uNW��%�aǊ
����g]!�~�
��9�-	I�[�E�OQ�N8}w�-�Fm4�j<7��.δ*.vA]i��(��3��a��[����tTux���������_�S��&�����*~1y4̦t�� <3�y�`3�����;�_c�j�F���͝4Ť�|~��[P��\�$Қ���P"���Tm=�qxW*mL����:�R��C���̟�yʏ[��冷Kh��}�(�9���X�H[�?�篅���k9��1����'Ç�CL$�^�M��
6�bp�<�� ok�A,6��PZ
K8�&7[�q��~�~`e��s݇ �q��:�(O8����/��N$��������������n{r%�����Ð
߻����"Z���^���7u'#��X����?�Ԃ��k�{檘�c=��![��`���!OG���5u�W���-�-�'��F�S�����t����}"�~��͜�`Es�̑���W>6:�wo~bA���9�>E��:�ϳ��jp2�_~��ꯒ������t}`G����]A_])��ޛ�P�SU0Q@���h�4�I(�9t W��K~�@G1�O<{h���T�^�Dl��#AI��R��?ݦ�[r�a=��?B�V��4O� ����%!�m+S9�~����s%����x�ʣ��*Uٯ�V�VF�l8ˎ��^!���By7�\�Kx���<Ų�>2�m�f�=�9��Q��������lEa��A	]����1̿���*4�I�+'�o��/y9n�h�t��k��ΰ���"�V���Q�XE��M�|��*���`Ĺ��/�D���cZM%�T�2�Y���*g�m	j'_�խ� ���>�=�brUu��������2��BcѼx�s�'�IK�g�ޘ�p��C6a&M:T 2����d��;<�L+�X�Y�0f���֧?�-�ϓ�tjj��:�@�bmX��X�=��P�Ѧ��+]:~���C#��������5E��h:���N̮�h�H��o jW����4o��&�TTss��p|^�;׏�z��*]蹉06y �l�_�:��h�X���{��<ɖ���-�~�P��w��؂��ߡ2S���͝D;7��U70�Z��B;�3�<�F�Irݏ�R,ui@���Y���^[�9ٵ��ך7����mLU-bA�����@��NQ��tt���o�5&��4��
�;���i;��|�,`��s� ������G�{Y=I�"b�1�ٞ��;!2�ȗ'��=��x��&T�1`��Q��,���a�|�8D��)ճC�Q7ִ\O�h�/�(�=�-�_jĨ�T�/���7\����2���(������\���
���v�Xh��J����%�6���e\4�ͷ�.S|]~���o��`��<.�<mG�����Ȍ���B5�VXT�t!B��Q@����ѹ��[�$��%O,R�'[|��)���IL�?�v U�� �<�ɛUi���Ĳ�<F����ɦ&���uQ"'�¤	���x�������ub�4t^/�-�ߚ�b{%nx�ى�<����1��2�>�]<Y�d��{�dGv�#�̵�m�|��T�1(|��R��+��}%�Z���֢�&������-�k��ճ����fr^��,TMzfWD�v���}w)�s��_�GNp��Y�_�"������%ɠ%�a/$�Yf��^GFӋ~ʳI�c�Ӊ��ڼF���5�%Z�"�Û�0��<"�Wj:�o���������<�C^rQzNh��-���ʶ��_`�fM�d��J����;$���w� u�M�z�.�%���d0�f��a+N4��G� u�Zl��s�l�|�l��9��%j>YN�������3l��M-�E�^���K�Jzt�� t�9�j� &����N4��+� ٳ�3{��;dP���Y���te��,�]���5)�C��Dm�Z7}O�!Jt�sÂ�H>DZgo�3Z���0����D(Ss >�g�i�U��8N��\�1��Nx�w�4��т�\ A,�I��i��V��� j0�>+;t��{f���T=�%�׻�'�%��b���(k��}x�t}�I)c��NC
͓1N�
�G���X�E���E�T(y�2�L�K�1��~�Z_\hH;��d��Z�]�Y�E��k���0CCH�y�K7D��bØ��e8,�,G��61� �*x��gx�#�T0k*�N3��	Oy"nF�z9,�;˟��}�#K��lCa�D�_C�+�ڗ��.�^㣠J�ks�vZ�;,�u>�G�^�=$k�B,��0��*;�f�T�M1e|�O�I��*�I`.M���)��ғ�R�U>Dyې�IL�G)0�hXƺw#b�a�*k
 �;���p�{I �QK�ǘܸ���(�2����v�X�V=K����y��{o���l8;߅��v���I�ò�����"[(2�G�w��1�yj�:�?���9���#�t�]e�\7��
w"��L��~�@��ME9]pif�h�x��^��y1���5�13�hh&w�>t-|г�bF �9�V"�#�q a�ڎ(��E|���aA^-�L�ʹ�̗�r<\���7�h��ۋ5%�P<��u~:��#%�V|�W,�s\b��1�$�Q4���'��B̴fF�6KÁ�X��C3������������{�=��+%�t��|�p�q���i�`<�D	@fV���������V㽟9-&�9�w�e+�J�l{g��1�^7!���Gv5Qt}�R [G��V�X�m"liS���y�:IF�=��+U��n��%y�{�J�A����p&��lP�+� ���بW��_�d�^�Qn_�R� �%����iT�e�{�6�Zf�4	�co�Ԧԥ�&�\87U�8�/��ޭ;d��ag*j�4��y��P��Y����.��8��9k��[@�F$�wԊ� ,SV\�Sg��Y����o��(ѯ�>�����T� ����Yj?~a%��I��hd���Z�<@\���f;s��t�$C�*&|�/�-~�4F8$�-�g:����9�سL?�Y</�~�������`�XXB�]yF'���Wל9#Py]�t?���͝hzVa^���9�q����97�����y�r����<��$�!�W����]�߿sR�v�<��Y7bQ0(�S�Bj���&�
 ([$�!H�<ރgJ���.�*�z�����vpKĞMF�:d��ۉ�܋#��}@��o���mMgFh@�_􁖹�R��u����maSN�(�T�SEξ��ŞN�y�� .]K�tpo�5�\OU�ke���AA�vS��[����������I'�������Dg|(ǐ��JU�ڿ�x�q%ضBW�x�3%H�m�%N�7[����k+�tJU[D)��M4W>y-Z�c����s�N&��WO�G�@/D����D*+�7X�..���+|�x��03VSxY����>��	Am2\-n�SuLI�Ir�I�4�us�*���j^�N�F'+�8AnyQU�(*�;��{�X60%�A[g~t���<!�Є�s��֍�:/�Q����XKY)w�p���f�Q�cN��}�H_x5�*���N53� 0{�)n>%��o6�jǇ1���W[�p��s3ß,1�V$�<>WNJ�8n��׀�!(iK7?����)�F5�$�{����b�|��ǃ~E�������B/	�9se�-?�ԡ���^�����y�g������u��]�p�5y�w/�ڌnKϡ#p�Q�=@�d6M���]4�ҿ�Z6E��58��&�-�(�ݵ�d1]�QH��>�6�Ȟx狾�*:�Ȏ
��28�7Yʳ�0��;|/%�S�:e���,�*�+���ҿ�6�.������NV�|"�Ŕ6e��ؔk��i�E���j��;]���;�	�ŕ.��e+
�lީ��2׀&��{�+�����+�(m�Q�i��U�%ݛj��b73@�;���P%*��WXX�

�[�︓U�Z0�f؉NB=��{��rL�\�9�XW����P�=������a޿IFv�+�](Uk�4%�����7ב��[]�����f�lSP%��9������P7�6��Ǎ�0�>�ȅٓd�{cX��A��<�OB��F��	B9��K�E����뇿B$k�$Lz95��ܽA�C�EO�U+�Y�2�Ӓ��	C��4#м]�5Ϟ�;g�0"S��X���jF3{ՠ��^s-�j3�}l���N�%y����\�Ne��{|�,�����z#"L4���	`���y��� ��2����v%�	K�pw�3�	�};�17�Јq�Զ�2��jO�������|N.y�Bz~���z�s_���>�#VL��?�����_w���{�J�R��A~��n��������V�0��w��Q����N�%�Z��j�P*���~���x{mF�C]��;P��(��r!I�DS�cSr@e3���q��ߐN�e����^��
\���O��)�%��A���\��=
ڭ�w�X�d�:��aK\B�{���-1�B�CeZ�h�=Q�뼵@�[HY�N~�#�ܑ
�J�LJ�[ݒ�h� :�Ia���o��*����8rd���0���D��O&� �����2t�R�w��0Rs*� ZZ�p�jRYa+�Gܭ�����h�,����l�r0D>e����Qa��J�T�L��G���pny-D���3K�]fQ�:������O�~�%:&_VNk�����W�&ӱ��3��&:� ����{��g����a���J��A@@���5�I�gw�|5�=S��7��®G�h����T��Է�YԀ�h�Z�t(R ��{�Q���W4�W��p���CCΜ<w�W�����
�~@�=:���X�%ʠ�I�B��]�spE!2G��z�`��ܔ�Wl�5�t��.�"����s���)���&�;r,�d��	�t:<^�B�Pi�֦��Nv�B�F���|�K^#��ۀP����~�-`��Ļ��e��/��Vc�(	�����>�{����1B����H��s���&_��V�F<|��y�����������I�?`�,�O��BI\j<�b�Mj<�3�'h�:+��+x-(1}�Dh�H'�@�Ѷ�07h	JyR��s�C���k	X�χ9h���p �^��&'`�������\��lM�?���[�$�5�F�RHO&�-`Oq՚֛Hs`�4U�Ϥm�_�e��|ٹ�v7ɜ^�� ��h�B]}Y`A9~7"��@	�m4�N�q��PE5�a�gU�w4�"�V�3R�v\Ia���3b�+y�U��E�����Q�(�,���z�i���q��ꉂeǻ��=UEKx5�����!	S�Y@��ˆ��I�xd�/4�����>�8���%SL��=��K�}�ʛH������б+%̸E<"�Li��~����c0:�6$*FoB��t��?�N�$3�Xn11$-����8���@v%�7VX:`�G�qJ��]����B���n�&(�W$�E�V�71�f~��ɤX��?�_��P�&��i�%���p�}#�Ӂ��r ԦҙP�6����QU>��	.�It8������-���T�[�Z�Cm��2%�V��M�FH���Q"��j���WZ���}�S�)�����)F�oCX�d<R�@�D�����(��,*�=$�Ҝ�~����n�uβ5]��/��N9���2L�����'QL��� 6�`���+bW�I���r1��V�~�e�}�dK;]2�P��4E���btG-)]�P���gG�6(\�'-)����\��D#��p��Fv������=�Ӆ���ڡ�XӪ%�kj��z�.~-�k!U��IS0���#�G+�ӎ����'��v��O�]��G��8˵`���bꪑ�p,4Ζ�weՂ1��=�*XjN=��_�3[B{5p��f��`����̲��n���8�i�����&����g��&�?f,6"���5]X��Q�]�}���)�-�N�8�0D9�@� ��Fm�0E�{�Y0��|=2�uNb
=�S��-�
���ҖV D\�T�ɀBݪ�^��V�ޓ�� B�P&���>�rj�}���6�	�Ex�K�؄�[�	���V+��fL����}�p�\�ҲB���WuR\1��}j����xТ;!r�qȒ�Qy�<��}�.vKD�!�qo(5p"	*��]��+ w'�b|ϩ>,����= +�]|v�ڬ�,@��ɀ�����V���\Q�Ϣ�c骾����Oa��pO�\+N��c�48�첢p�����q�3DO�k��Ԋ�^�e$���h9no�l��M/-���A#���0$;M��i֙��X��|�%d:p)�y�=z}m&_N��(�a�Ut���MЕ�p��/����	d�
(��[6W`��6�*f1�0"81��P�.j{��EÂ˾ "�f���q�6�����!�s�OD���dI(��Ƕ�Yy�ә=4�s�莏]��K��/��Ob8����k�-���ɸr�rh	ңl�����|���7���m�e>O�����= 6@]�ῢ�S\��d%ˀ�_���?��3�~���JxnAE��P�R�~���sC����<�3[����[����D'���l�U.�PQ�7�m����،�^��1H���}��Q<�Ro#/m9و:8���ס�s"���mGբ.�^���s8뢵e� �#rwe�:2}�P�L���ڌR4޼���2�����S���H�f9x"~�' ���h{D��R���W�����C�!��K��JԜ��s�ς��o�<�"�K�!i	Q�5�~PR�G�f�g�_�OH��M�\�����$�ESdٞ��������A��90����8a�2�H���0���9Ż��6��A����?[(>/16�ZKy��<��]6��z��>nYp�g�0��f�B(Iђ�`�2Z���RnIf:�d����^ۂI�+���}K�qP�_�� 3�S�I�\�o�����q1Ֆzz��wNː\�AO�����˹�l��0LS�2��ڠ�H�*�juw2=�9��c+�^�&ʊ��;���ce����n��c٢���	ԧ'��n�9��H/ｒ?�,a�c��Y�?iL��~gY������ҳ����D�yHo��@�J�
����tm[-(O�S;���+k����W��"�|"���$_��q>0�%�y������s|��B� ��(_7@��B+Xz9��Y� �?��Ĭ����4��TO�������*��R.Mg�Y�|e�����fआy!�fM���w��+9N�I$ۚ͑N�~i�0���Yȼ��P�/��t��<�f�X�9��7��Vݑ���J?M��"�������p<L�A,W
��۰� s�sF�nǆnZ*v���ė�BP=�@�:���!7*fz���zVĔ�d~@4r�[/f|�������b>�T�qfp+s���=!/>d��Ao��5o�8�~zL���샇7�ATf+b��J6�Np.*����)o���U@�e�ͯjP �?�Y �C��J�0��gF�g|ur��/ɦ��y��C2-�(+Xq6��;j�~���	��O� `G��<
nWH��R��G�޷Do�s��OE�/�M���9�a��VW�:����}���6/h��a�,W�d6��Wn�T���<B��E�2-�M'&�� $�d0���c���rz�d_�B7ݫ�<�'a�ي^�9�@\�Ji|���(&���9c��nz��
:�̈́^��M��Nz��VBw"m�"ٗB�j� [�`9�`xdBՖ����z��}�����;:��n�R��q���/E|��S��\25F���#|D|�.�e��⃐�Y�|6��1�Q7t�����CRiV������/}XA�jC����a4!��]�CEs��:�y���e��/�}�?Vq8�I� 3,��^F�e%_NE��r��;J�:�n�ħ�_Kb��~���E>h��{s~L,9��Y{a���ￊvЛ²*��Ƅ��hٯ:&�ו
�D�Y^����j�u�����RyO�C~[9�O�m=�a+�IymOJ��K�y0���r�H᫜���1+��������!�n�YA���j��I���>M�+D/5���ط�I����Ց����=޸��b��%I�e�HP��`�hq�h�>��"�����%��FW��,�4�'G�۰	��q���
��J�~��x��3��+�6�^Qˏ�#����vB��|���υDs���e����RVa\~��hJZ���y@�`���Uz
�{/8}�2�ko8ko�c'\{��k��4�U!6���و��j>�c&�=6������]����h�R���+�� ���7�bJ��QobO��B]�YM5b ?5�;������ܔ�\aB���,��Ht$��5���1�����ET�"����{�M��k���߽�t�j��sv�[�����Kq�i�H��;�R�bWz���څd��3�mGh�$����ji�� $N�պ.��I�s��!�Ҍ`0�X	�Cf{�]A)��ίYN��@���I�6�MZu&"<�b��qz^���4�m]�	��ez��j��d#�z�ܤB�&��e�d_v��[D�jjdmρ�젆�T\}��Vz��Nk��G��C/4Zw�F�%R/u.��D%�� ��������9�#�Í����5%ͮ`a���A��7��u�&��J�(�Sk�}`Ό��|�����I�s��Sczr�4�c�����O�B]���ڞ���&I����hR�؜��Y.Y%Q���:���)l�,;䃳�MY���rY�s�\/6��YP��r�gk65�m��M���U�o���E}tvs(M�0�6�nj��c e�HB� IW�7�s�h�8N�`.�O��a��Od7�#+�b���<ƶ��Tr�sT��e(���������}�_��Ҫ�Бp<���}2�6��ɡ��K��K\ɵ=��⵷hG�
#OmY�~�D�ǩ����c>� 设��,S=�S��Aޑmɩ�6H!�s���	�%�u�^�q����+�{ZP^<	�8��¹�H�ɡI�v3�?�7Wœn��
`�6� B١o���ї���Q3N?�q|�Pa�a A~��p�]�Щų���2V^}�:�	?P�Gf��f�p�M���e�vm[�m�h������|�k�T����+��\������E��'����)@,���T��\�Ex�@��Y��^ܶ �"��N����rY]��W�p���=�fX�訡$PE�2�4���y����-cmV�3�$Hm��f����|����;����~&{�A0�a��tp��e݋������'-���Ѡte=�7�s��I \7��p�2 �r �x��ീ�
�jm�A��$�_F<v���I�cȐ���Ǣ�kMe�� y2�A��\J���<��-)����[�"����)fc&3�mcK�%�\�*DAk9ybX����eY�b��ب�Qp�8�Xl@�r���͸<�ͣ}v���'��0pb�9̲dXO9��.��==��B�|���k��(�^��ZI/}2���y��5��G��I��DgRr�jNͻ\ a[gB(�Ju�x?*פ������s��Vy\y��lɹ�4ٙ�џ{bT�r�:��S�B�7$��&K��̞�DVe�=�/�ِ�4���U ��ְ:6��f�- U�۬�	┹���p��_i����g�'��Q��m$��&K�5�!�;���/%FF��j	]g�C�{&"`%���P���E��Ҍs��9�hR�Ʃ�w}�/|�Z���I����?2S�b�]G��7��\�_�� ȣ���9{�a&ք���2�>��~��x��<Q0��s����QId_"y}UK��{�y�]�3���/����]_2�J�^�dp�y�1@M1�8��*#�Y����.i�۱�[1��@�I�e�a�׿��9���p�h�YS�[u��I 5�JH��3��_�8����dӨ;;Snu��{��W��F�ŪJ�~�o>1�qyb`|�e�ٯq3�Q�g��j��gcJ�M|/��`�Q�L��hbť!���j�Ȳ/�I������� ⿳Fe��}��a�J���47�᫞.��,�
Pfk����G=�N��d9�ظ���[5��S�JK*���ƶ��\��S��P��/�l|���ӈ]R���	�*b���t�K^��`C�?��9y�� "����J��A5�r-Ń���\l��GuѼ��nd�v�ۜ��c��`�h�c�&š�g݀@caP/����'���6��V��n��\>���<o�ƞ6�_`J)�9�tc��݈���_$� у�\�"b��ִΟF���`��>�e�َ8j������ݢHDa�v�[z�T��tJ�}���Ν�_�S��lD �T���k�+SpD,��dvo���D$��-^�ܭ̈́!!��:Y7Ep�w��.���:����:�qG�З�QX¹�l��C-�<W�sʈ9M྿��%���k,�9 �]��'-�1�+2<8Xǀ�P͌׵Z䑍��z�p��n�@��	P��t�)/�[�X�E�<��UָW����������ܐ������H4;9�P+���+,1�	x�~F�	 ��&x��f�ۣ}����F��̋C�)�$�Z3j𻖔~���"m�� �L�pO,o�&����@}��G�Q�������l��E�T�H�-5�n9����{6��l����=lq��k(��{@3
ˮ���>�\��vQJi�o^Hځ��%�W@�ٷ��u���[���̪��I��(#��~�������~_��wZ^���y�ɜ��#�A�ߍ�s4�c��g�.��	w��|� �E�2�Î�U�%D<X��������&�Ƴ=�{� ��ڻZ�v2�;I�_�'_���E7cx��p&@_��(�_�X�|)�:�N�<�O�m��6�E1��!hF����Z���=����l�?�J�oY�����\#M�x�xȢ�=�����_�kI�`75n&��M�T;HO�CPx;μ,��:z��m�������ɿ\�� �_��.@�]�FtgN�i���Z({pZ��#H�`�L�s����ǤI��)jE��}�ξ����%'	FJ�Ƥ�!�[�jr�t�)|��h3d���F�*�#w���RQm�7���c$l��v�~�=��|���ۨ��2���=��lI�%�.�n &�n�9ȑY���ߕ�r�]>4��U��;���|Eo�� �jH�Z���u�W~�=����g|Ae�l>}ڢe��(ήi.�;_��2b�i�����3�7��a�Y��Y�**ѹ6]e�!T���OF������gV��c��~��Is�6�繓������W#p�'��`�t�����V�#RVc�.j)�<~�(�,ÈE�a6�W����.7���>vlz��Y���Bpl5
��1����T+k9��y�\3�oD,�n��?dv�]-(����M�m�U�#���d�Еx9Y��`vI�y�cP�PPȦ�j;dcE�����9�L�Z�#!
����v���T���Ku���y�ω���{P�3��<�&j�x*�q�mh;P�Y_~�mHz���Z$\'�:��N�o�E�B�yA0�`j]��c� �3�� _bP
�����%x]�f*�-�h_h��7�_9G��
�V���\��m>��zݩ�|��?�,�ӓ�y��bi�E�ϙF^oGKI8R����-�?o%�H4/v�\��vxִ�l���W�w�1�C��˙�=�)��l^�T*C/�0|\�i]���Du��zj1
���Wt�S'R� �~3FA $��x�BՔ��3�C����������ͥ	�>[�1�۹�|R���v���pX��0��z�T/��c�B�f�P�k�W���S�,��N�Q��77�kU�w/�d4���S�.���5��yy�G�ȋe�D36���A�菳�����#Q�u����M��!p��<�ޮ�D�;[w�lsX�<l¸x���q���J;�l1Dޡ,u_�tS��"�n����cD�4|,��=P�j��T��s�2r���?!�=�9iPW�]7�9V���R��5F����`�b��f�C\���!��_�������b��)ez'�o*�?��m�������<��9&3��?�`W~[���I�jL��_�s`|��V���/M�{�z�<D�&�_��?(�^Ę(����hj[P	�<k�����C�����P���I��5gyxI��k#�o�
���a���?-�ɸ����^�Q�� !���n��f�i�k�S��kRv�o�KW<�2����	��o��N�l֞��

�P�8&��ܚ�t�(����gw짩���wQ����7�a�6c�~UP2���CY!�8o�l:)f��>�'�],����J����.1�ޯ��<�q��`l�N|��H��=��� �%Z1��z/ě�dJY2� ~6�p���_� 2�4�L)k��y��E�`��\���h`����r:�d��e��q{�ߘ�#Z��b��n�b=ހ�A��8��B 9��B�tw���#���D�U&��˸�����|��&�cȢ��џ��7X������y�.�P�ՓS�-�\�E�݄��R�@E�E�3���L�>��Y�YB��SZ1]��1�PH��ӄ�����m_U�^�۟�`;��mwe��{��X�f�^Z�t)�n�ү��o ��m�A���[jF�+2'����/������˻�eX~���>�qG��L�^2�>:�6�e-�Ü���۵Ex=���>���|��*�<2���Cfш�'R��U���y��(����iZ���"���>���Ӌ/���%:0��'�Y�<�~�O��Pj���&�����&V�Q&�\`c��
�%Dg^�A�t/̃�b|��#y��5� �B�k>����a_\I�D�K33+��6�)�צ&�V��%����Ė`���e�1b+�h*>E+�f���z+�Ds0BK7w?R�ۙr�)��w	��H���].�j]"�]եg�%�6���)!~F�?��O�w�U��g�ެ,H�	���J��I7`�r������
'���W'�a��Qo
A
����t���o{�|['m���t�qk����)�U7~*^W��H�?ßF�Q�9�z}(gk��Z����Բf�����_E2F�{`��x����z=��᪙�����T��G���ƽ��M�m�0�q��v�-��<�݄v&���̸����=�#RY�%Ck�D
����4*��I�aL{𴅺�\t��ߴO�EUM|E�r�Fp��(<�S��N�p�����M�[�����XŦѽ�Q��q��o��}�T�ΆӥjZ�	08y?�0�iorB��j$9j�qЀb�B0����Z���3�|zW} ��p���}RYTFs��U�
Tin2�O��S����ioIO#��=�y�Q�k���Z_�n@��i��CTM��g
��'$A��`����NV*���;��  [ �H����Y��8�^��z��(o�H��bP_/ϴ��=���ܤM{2�/��dnL)̢�֓[���Œ���d:4�sT�kuS�0��8j�֭&`���D$��D�V�k��OzO \_|`��B���h���G�-b^�g��Q�Q�.�؆�@7|�hF��n����5S��~D����^5�1�y�����'��Ι�=̗��@"���LfW�Tv4��?��a�1+����vi�y:��'cs���&���1`��O)FfF�����iA�l\�>a�Tk���]�uې �?h��B�h��"�Wp�p<�-N����v�f��C�G�����sh��{)��1
vׯ�[�åq[tOM��	��K�e�m}��j�J�e �o��#N��
��1���~��<,[���p�2������� k�����!FӍ~��(��o��}��<E>jJs"Q�PnK�� ����F�%b�J��8�e[n����`B�d��˄�r����o>/!.ui�Z�y��ʙ膪_��F8B�\D�����YR�S�K�3��V��S�8�+�_Y����ۋ���v��(��H,���qV�"��\az�'�goK�V|�8���W5O�B��/=�:2�m������l���=�C��3@g"Q��| ??��8��}��+�� ʫ	܁������/�v[m%.���,�-�iT��l���!�%O¡�=���Rλ���z���lp;7�-���ny^G�1�{;N� �o[��G��4��¯ɥ��5�v!nl���l�C�ijϣ�lV�G��i���c]�8�����a�N1V�P#�鬚�E2�C`�t$
� y!�\Ç��r:jZ������p"����v�#I�q���:�{� ��'��0�lH�� 1�3��W�D�L����??V�%;�q�u��l!���~�����QI-�Y�D��z����#ƫ\	�iR��x`ı���� :��k��-jP���&'EP��;-��/0=.�5��+���K��\՛��џs�
ۚУ�؜�1����u [|���}j��g�K�ٗ��42ee=�:zԕ��$�g(L�o,~rJ�'W`����Z��4F�4�N�S`>�L^���Egς3������o^}�6�X��AS�j��23�.�Io����0�M�