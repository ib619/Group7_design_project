��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����Y_��F��tw�p�^�=�����DW!of�.��"�"V�8��Ua}W#R�M�-Q�xq��ų�����#k_Q��?���B8I��c��l��{ͪNȽ�D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����~�Yp�Ƹ9k��*����l���˩��s�u#���x�} �^�<�괠�<����� -Ч�<3,6����*�?:���R���yK�q`Ĳ0�Bܻ�����Z\ʔ��+��mk̈́|��'DY������n�����b7~tr�cm��נ�U6�7�sP�����ߏ"L�H�,j���-\+��W�ā�(��7-�+b���46��8B��16��'��~�C�u��{���0�w�C�rZ�=�Ft #�`Q�����o^� �L�����nY3;�'*���_I�淨Y.އz��w�6�mIKx_��S�8Ḕضݝ?��RD�H�k6�_�=kG}��H�15u�Ԭ�����)>t�b�zIf�6���3`Ł��#�o,1���mn3��/_	�Ѝa�hg�7�/$�:C�`&���`)Y�^�Q߫�ޭ�hQV��2?����X�Ӧ���9�S�i��3����h��Z����W<;����訧/\zZ�����^��$X�^f�(�Ŵ�ā�孏[�L�@��vۻC��!���F���m�mڵ�k}X<2Lx�ϼ�o>��g&-�m��[iٯ��w�m��	Cé�~l1 -�J�i<F4���l�/s�"l�;F�Y�M
�\0�Z��e�~\���o���ٿK�H�|q}�iz�K�K��6u�2KE��r!��Y�Fm�W�&^�����ޘźMʃ�ɨn�C�B�����%~� �ӻ�13�J	���_O��B2#�S8n)�K����8�No�I$ ��Wy��� ��@f��p�z�Zu�8��<�b�e?�b��7r=�0����g�u�RQw|Q������F(ɓL��5˭�����/"\*���ȯ�m:���N��K��'�_�̅����#���;�˘�1��7 �iv"�qUg�8�F^�����b���D�I�*7�Ո�N�ݦwQ�ȿ�Wͪp������rP����jS|$�w0M!&icoۻ�>'a_l�`Y_L������j��UN�=�_��`!�~6f�o�Y`)�����;5+?��ջ�z�nP��D��h���2�a��ۆPKa���jg��bc��a��<%����z���bk��\K!e@'G�µ�̝�
R+F����a�xcU!e�����7� c��L�D�(��\�,m��(�o7y+��5����>��A�2`�q�����B��Z]�t7G��
3X�?	h+���Ka��ŏ�o%~��юz)���k�\�+%^��%"�ef���ج����&4��UX��p��	c((%���xt_��Thk��ڷkV������bQ� `ԑZ/�ǋjև��5!���<�H��3/����V:��z�i�#�T�K�ܐ&����/�R/^���~���<g����o�SU=��ϥ�r�t|oV�����G�o�Vl19�����'p�ХjE���8=�DY��E.�]0���G�4�Ik�R��F���o��Uu��:�%�b1ݎs�2x<Ż�H�?�Aɇ��s������a�	���\�� x���A��3ȠQ\!#��E� ;g`�:ȼy��3�1����{�x�����{S8��H����i�`�k�5�(_�$��BG8���F�CJ׮!JRy��xI2뱢�£S���҇��Y!���&�|��.>`n�T��y��@#�� ��]i�.`�|�Lp_W���#|��$Z��%�;Z:L�-�ϵ%�9UjcuM-���}���79'1���ׅ<6�?&�7�,�Р~�9���ޥ�A����5��*��"U��W������"Փ�NI:���e ,y�q!\��^�)>��r�p~��V��-��Y���(a�Aw
�����V}�nCt����e�3�r����6�PX}��JN5�3�>�}�
>�CO���Ҙ^, zv$d�r)�Gf�#@��!�(h����ǖ�Ӳ�G�� �2?��RL$����e���� q�K���8��\���z2X��7,�[>ob�q'uaw+�рM'��.��[F�����O����R8�}�*��(<\��f��b��[�8��c�/��#KV~;��`� ��|kA�&w����)�H��1�B8�P����:���*D�ѯ�������A�=F3�_$���ҁ�Ͻx��A����� 8�{i+62%:�ڦm�Of|x�#'��ۅ�-���d/n�q=��'E��!��+)�o�U�(�|�f�ޡ�e.��V�ŪG
�,��	������ܠCL�B���[1�C��:˸�ԶT�,
&��{`-����VI"����2�̃q�Dg������g�y˒� ���U���;c�w&+��3��*N������`D-��3!���=#�w�P��C�KhK�tF� �ڹ��y ��>k��짹ϊ9�E����'L0�-�E�ƈ��Z�b�!�DV���V����Z�
��I�"5t�e�� �j��n|�۝�}5��gޖJe�[ro������	Ǯ
QMx��Iс�=�FS�|>�}���H�-�����#�E�H��H����Ub�xo�bH���F�:�������$6�b �W�s2��Hԋ���ⳇ逶�۠�k�/W<�q���y�â����@bis�%?f}�|A��E�*�?^�N���Te����n��6_jr�x��l�N~X7�>�I,Ի����C1���-\����@�����.\#�7�]�&�|ڈ�ɚ\�|����j�5�~���ldx랃�j�r�"D��)����~d^��zj+-��y��	�˲�d�z�p?:�p�$W��X�bv��kW>������`'勼��_�t�@������L;~ݍ����Ԟt�j�E���յE�|'��VK�	ޔ�"|LY�u�����U���1�.�� �brm:DR^�
 zP�z#y/Z����(tq��QN�0D�����@Ť�fLD�w$�[Ҝ��o}m;�����z9��,Ulxy�q�)����1���0�ê�1�иp-���uT���Lm�8����B�+��	F8���v��R���C
�&~�K���4r��:���e��7#��!j�UY!.�3Ձ���6�BQ�������M2���4�w'�'��d�s]����jb3���e/�56�z�2`漻W�D#�������JVȦ#2M��F[ ~u��V�g����d��W������E�����g�Q�=Tl�c�~��,�<���E�*ϵ��-®�}u������:��8�e��V������0����(�{c^۵0D���0��Qo���=�ks)��e�|v�^��m�3��g�؄�&���j���K.��Ɏ���ש6��ؽ�A7�^�r�t�m�ң �L>d	�����FĞ�9��0��?�w����ŭ��j�"�0u�884c�JˉE\Fƍ>"T�A�jJM��)ׅd�OU��Q	�b��Zy� r� �_�,$��0���=�y��(���ۏr���*��XK���ܕyA�E`%.P$,|�E���U�p�����m3D�_9t�zc�������EMI��M��ޒ����nh�`���5+�X�O{�f��p����.�<Y������NF��;"=��� 5����>	�HA�_�.�s0ܵ��!��mr�䆲��4	���J�qA��d1̱�Q���'�]��h1#D����Ss��df�+B��e����NІ����P"�[��9N\7U�ޯ�]1@�T���.[t����-В�0q\���S����1�o�����i�s�P|"������t����ͳ�B�z��1�:&!җ� )ȧ��瞥H?!Ѹ�֌�I�i�ʐUqN��!�RED���f9^�鿗�Ay�)���c�H\6��l�A
;��ݻ����a *�F��ܝB4�]�Hf��I�Yc2��#���(�g�=�A�#}�m~(��'��?5� k�8�� �jO����J��9��E�����A5�I[�����UB�HN1�#���<B��+9Ji�E�h���ߒ�iO��տ����Q���L���t96��e�ܛM�����I���'�_���4���0�ϻ��������}4>�ʖi��mj!ɪ�H���H�����U��oT�~��'L���cə7F��8"on�E?L
�һ�d�#I/Uc�VHM<[�Q].�����\>?�wQ�k���C��d�ik��z���j��]�xAuYƘ�UՓ��	p��呖�Bk�̦����uԐ��J�}� �k6�s����s�;B�,⺊���=a���g���;&��Y� ���B��x��O`�>d��쬠�j&(��80'"!II�G._��1|��
��8�)f�Jp(�U/�A�M0�wO��J�E�C>� UU	���>�qLg-��}�Ou$p�ek�$Fea8�>GNd���T��o�R�� ��A�~°J-<���S|�MCKG���CC��w�܈'�;�|l�?Z\]�ֆI3����`3T�O���0���9P��Q��铴TM���Oн�5ޠX	Θh6��锛�(�un�H5�U�w�$��u�S��p"�rB�+aWBq(�_O�WQk������^��0������ޟ)���">�;�ߣ��eں�p�6��\+�E��8�����c3�T�e(.��A��A��="zy�%	q��Äf������$o7�o�'F����qw�.���R�vA�ΦA1��� ��������-�ع2�0+/�M��'h��G�]+�Y���{�u�g���`�"��,��4����7zL����=�@ �$��A����v=�m�R\���U��=k+f�����pOF��I���9ϽKH�E�u�@�A�ζw���va;� �b7��Aזi#'���bĺ���YoƆ+����Z2d\��d�Meƒ%�L��/���0�]3��Ԓ��[լ�b{d����9���N��K2F|����|����d��<r<�2��V2���j/,����ʃ�"(x��$W'��V��x����$�ǎ��0��5fn:���@����m�����J�["��I�W�J���sо:#GO��߄�7��1�(��)S�cGE��O)�˫��Hٱ�aw�8+���SRV�M�|�	�q�(��\�VC؊ޢJ�#�Ӷ+��K4��1�z������Z�о�|s-.��>��|��1%�N��]��=>0\k^Yo(��I�([h^'�Z���[�C�c�W���c^la��U����.zu�g7�|<���ӌ��g��w����t��X~�x������u7%>���V9��ѝ�vˤ�#�ww�$C9�`�D����ߣ��d1���p�t,ù�I������(�<ћt���A�ajؓ#7e��P�������N0�3 K{����g%��AD��Vl �7��K����M{�6?<(�}45����5.Q����*���%����1+Xh�`�h X�����0�O���jmD���H����%��Z�J����'�`OS?���& �3I@��|i���<A$(���������DH�|aN�z1��˟}�W� ����Q��	��U�#�����;�*�:��ԂN��_�G��ol`���`D�X�[m��L綔���Q����հP��o�g��H�E^�'hAp��@��߇|��b� ~�e7+��+�.��3�nT/0���#X2YM's�47�DF-+ys �g��S�������f��1���7����,>� $�ÑY�)$��8�eL��p��X���_���6ΗNr"�u��-�����^�����Ӕ��5�z�<�,����F�[a1���n��I�}rV��/@7[R��u���D�\�����m�eފ^�N2<Z-�O��+�x�"5�
h����RV�UZ��n�#m����R}��<��v�5�*���Q�L!����r�\L�2KI+6qlk�ϓ���&~RB�:	%�"�X}�tyU����3���>O�(�f��!�@�S�����v�~ <D��h�Wp�Lb�(t������qr)t����[Dn��?����1=�#��z`�����?J<����פ���R�ڥ�:�f�>S�v�|
����ʛ�QfTѱ�\�:T�6I+s�on@~N�Ԛp����w���%[��KgJcH�Q�ф�MW�+"���W���u����vT� #�Ĕq�C�؄w��Hk�Y���P,Es��P�8�&D`�����O��9���T,<�H��AF����p�Iٲ�â�h�^Eo��=�X�`>�z��ŵ+U�[�S֌��:��Ö�o�~��O�B���G�R�e�cgi�d��o�!]�����q]��y���`o8��Pm:��t�j4��4�����_��wp֤�"�H�+�,h������#}<ꃔ�=9˸w���ed�R�GP�%F�6s����Ya�Ȗ������Q�����u��ZхȽz6�n���د�ݯw�iL�d������dg�zAb]�]B�P��ϥH/�z�Krr�?��oc08O��PՀ�̚	5����r����5�����
v�ÓL��}P
���s���4S ,��h1s��/�������S�e?f�> �M������,�lz��K�#�t������_�
�8:9�<)Zf�$�cb��C��~�����^vߦ�>M�)�ƝZ���7�_�2�x�ݳ��� ��ŗ�B�a�4Qd3�%��R�H>&��y�����3^VCu]�1�m�Yį�*u�Q�ѷsغ,Ѩ���)i��^��wX�O�G�5f�N��~����C�7��6xah���]Q�w@�n�����4�K�ǎ`��&�#�2����#u�R������hE4�A��l��纅A�`56��$!l��i�l^�	��T���fZ؎;.C�8��
D�jm�H���
k�E* H�b&��̥jIb�lWro�ӷ
�"YC��,�CC2Z�N`�������V��ĥ�~�Sw����¸m�B����	�1i&mHO?3��N(?�8��@��r�b)�Q����Z�~u���ܜ�?�F�Q�Z6^�]|o�x�Y�O�>���t q^���W~���}�Ig���W�/l����V�[�֎S쨜�{��*�T�h�U�����=�p�u���l���_�lw��8o�Փl���%��NDd��P�d��ߖ��ƩM��􄒉�[�U� 6̿\Y�W���3e?�Z�9�`�m-u!s!4���q��8���6e�=��E��C�_Z~�\��e�\@�q���h�fa~�-����>A7=�WX�� �ArlU��������n�@0��S����E�o��,  :��D��0n���;���c�DX
w��0��73���1)�l��|a'?JGUWmpj��u`<���:Yp��&�f���uȻ\6H��6e�O����q6�����+���J��|P�0���kr�M��Vq�V7h�1Ax���W��5h �ܿ�K�$�Q�S�`�8؍u ������0��t�͡~�l����=����WҬT_���ꇰ%�,�>��f�o�/ ?��\K�hUbvK)S��w�D(��Ew6:Mr����.���y�9_�ʸ/NӑOm�;���-��j�T������%a��� s�T-$$�Yf��Eax0WW-�Ӫ`�)\�wN��<T�k�I�g}�eF1ǹ�s�\����P���3�g�ŃR�jrAt�ٙE����!��C������NV��)���K��ؔA��pY'�xvf>��Ů��>��ll��5Pp��ݱ�x[K��~�R5Ͻ���m٘��%t�^c$��o5��߃�G
{j�,���7Y~����xX0�lu.��
](�u��
��@ʅ��eXi9�!��c�4d3�����b�!�i�X��*Z�9�Pވ�l��*$i�B��� љ��Ђg7Or8����)��Ȥ=�Y��� .I�t�+�<�?�"�`QKdoE���'Z7 �=8��1�h��£4PE��#�.T�7�EB�{;��%���V���:H˵���c�L�x����frQ�i�P���A�zY�����:�^�7��:��ҽ ��Z~ݱX��`����f����0�8Ka0�Dq�</,b��D}7_s�塤�/݉He�ulFx�f���j�c����Ԝ��ok�g� �剒�]Ľ��KP�rk02���w@��Ny �v�ZMZ���P�cM�mߡ��� \�)єm��e�n����j�>Nw�������G3��O���rݙ�E���㌾�$� U�YՌ���6�cFn?�( v���^�*�s��E�����cN𕃧�iq�u_>�=J#��p�f_�ӭ!RJUpݬ���y���#�KDCO�ԭ�R~�]H��@T�TƖ���X�'��?�Z�l��O}��W�:��;�z����\���g
� l1�ކ/��ߐcr�S�t1���G�����h�qW���%~�=x��Ջ�
e>����,��A�՝��Lw"��}��
�*/��x��;WK�]�*�7������G��?l��F��/_�V��Z,����5��gЖ��$�2���~('Ro����Ϗ�Q���⾉�=�]W��d�05D�� :5�*�'i���.�9�a'$} �zo��͑�R-����:�<�uP8N
�य~d�!�=����P��/+UZ&#�� ���c�!OX��a�Ip��zS����V��V���a�s.��##�������<~p��M�{��1�LKi�u�3����?whUl£�Q�;�s1�6I#��	+�;�MBLSW֨~SW�|vĦ����S�������TҀ�����dܽ�$ MZjq!�*�#3�~�+��C]�OD�A��Z��#� ��q �'�Z>��rE�E��=򘈕 ;}ha*���=han]�D����K`�:���_w��<-o���/�[~sZ�m��ΩV�\t/*��A3��~��Wi���}�@�����F1"h����b]"^�oK�@s(�{�A�ߘ)`dYtzA�!�q�E�hc+��>jn� ù����J����G�"��Z~�GWR�fE �UmBA�5:��}X��P	�:V�|���� ��mXU��`�Ǒ_*�.�U�Ăl�\���QA��^尃�$�ܩ�ҥ6s(�7ɩmP�g�b���7k��H}Y���	�@���M���%4vP�Ѹ�V"���~�X��q�;DGܖS��a���q�[X�p+=�9�4�l��^T7(�'�F�*l��X:��(���y@y��[	 �#�����"ߞ���ym>�&t�F�Ng���M�|ܐf��~��%2|���W���X��~zqQ"��l��C#z�&��_�f�z. ���[l���)�➷�[մ9�{�E$ތ1_K��,�n�qӫ�:���)�;���H�%���ܚ����g���9'�#+�#`��e -�>�R#�ҋ5u���T:��8��,M��n���K�( �eы�tb��z����,����<V��n�c�R���t�\��G������Sūv��޲ڧ�@�tkT�=���[.[���:,��KAm�T���
e쌽/�f4M9L�#���*13 0	�ۗ^G�UY�x�P���r�Yd!��
I�2'v�;at [����(�h� ʪ�>B�usE��b܌mks��s�;�G]��з�8�L����)��˫�!�U���w�i�h�[��G �/����f�H&"�����)�ժW���ߝm�j��&Gc�9����0O��-�$����V������d SA�1~���WR�O�J۳����$�����!�Tug��z��]m?�ϖL��[#���6����p=��{c����:��`����n��ު�'U��z[��
�S~�SAj��Щ�W�@��������]�.��*���;���gM�p���2�F�.�A�?�d�&�����0��2�B�������鎌��e�����r�5@�#9��Y�>�M��Ѱ/|��:q��!E&�!�	G�Ӧ\���)A� �
���	� �|��~�Y$j�1R��֜n�B8�	X'�x$�����cH��U�K/�)�!�hxi���ʥ�%��j�L6�)��Y�y'�=hQ�\fJWe|�����a��2��Z��W�5���~�F�#��
�s���:���IC	ON��q�Z���[3s  Uv��08�F��)eb��C*� �g'���L'L�B�0M�� �[�@M���y�Q +j�����<SC�@�8+��;�ˆ�d�%/\�kwj��X�X����^gb��X���K�c ������|ZҎ�(R�l�L�ZNWDmM��`���\,X�%a���5�Y��G"�U+f�"U֟�� �}��%�6�*��'J�-���S!"
(Ĕ����Ko_��Z?��/ȑX4�g�o��2��NR��{tY
���~�O��FjE�,��fz��:;�7�<_��b�+�%�`p`�3u!�vv�p��u ��܀G�'J4	��G��J�ē�(f�㯯�Ǎ�Z�0ZX,8�=�W�q�b��ӞK����Ŭ�T�ͭn�M=����	����$�vK�{�MB������ᑣ�pпōce���S�+[�L9|y���$v��>PG@��nN����0����L�;h5�Jۗ4�A.kyj½K��$��v<��r��bL�"!��r�W��� ��$�7�akσ\��+-NA��@��-�p�emސi;��{Lv���8}�iW,E�t�ԅ����bN"Dj������7��;�V����Ks�֝���������]���Mt٥B�9��5-��ģk��13�'�I_�h�S�`h�>+$Gح�u@���n�Gj>
�@���V��/0[��7�J�<b|+)���J_�>�E/i��v����@R�>���H�o�&u�0��85��w�z�_����.dh�e؎�a���g�-����"��n�Y�Ĉ�y_�����Yb���n�wJM�R�_ĥ
$ۺN01]�Լ���B��?�F2���_��$T��d�X�\�����1��P+�tW�GƜ�a����nN�q%Jô���c����I�Sm��Mb�����g�'}��rRm��x��m�-�J�AV���<��u@Q�X5�?�b�r�w+)�����;؅�s�U��?x�ݷ�N$lS�!.�7�0.�;�]��n���sJ��K]ç��̜�g�ٌ�J<���қ�����V�,-i_Nd��\uˌLto�4/T�y�UT��Ȥ�*�QkǍ�6S*����H*^��n�F�rH��#���`�𗳐Ju�[������ wV�o�2��( �`�E2��
���u0��_k�k�1�"+���\fK����>X�ʷ�y����淲�#1��:��oe�?��_�M����!�=%T:n�~�{ O��&5'���FH���x�1Z���ɖ�b�������惱pWŋa�h��ؿ����.�Sgs���y0�F��kZ��l�9c+�y��\S̸��J������u�~8y�C��K��eJ9�x�*��>傳��2u뵩"n�LjF�@3�&�Q�#K������`��\����B����^�*��Ԗ�K$���Z7	���y}����}�59�0>�6}]2�U{������T����Iwn����]�)�$*��UA��}�ǈ��:�-��t��= ��F84ɑ��h�%$b�\NX��h|�J����b�,�L���t�'�5�D��\��?��>\P/�w�R�t�c�7�SY��~Y�4 6V���׭Ҥ`�<?�S����\�jNW��E��A��i�?����e`|S���))��
�a�~xD���c���kͨ�.͓;
3+ɑ�r
�K`��[�
��Ri�˰=�J2�����[�����\���q�� )�k�_�A9�G���6�>��Vs���q0
+7ȵ�t�G�@6�?���R��sdU?���C�z�c.�y5� ��6�=#���|' �O'+!�w�RT4ij�lQ��r��G!̚���jI�s=����S/���>l��ai�����h�\��PǍ,?�Γ[V� ��z5��>�He�$6w�[��Psf�#t�������=����vu��pc�g�����|�@���D�PN�j,J����o�T�j;�S�Y!��n_�D�
�
�c�2���":��G#���h�������9i�5�)�����-��?��g��n��W��0� /?�C��WY���eg�9e��Y�u&�p�����?v�d���߻=:�����H]P�WJr=��EbJ�V�i�r�pwpN�"��Ҏg����a��2%H_� kB�Rl�L��g�c�"��U���a�?����y�\���pa���|"�_q}�0��d��J�܇��s�Et��c�Fn�5�	���������U����|hH�EC��a�p9��Ʉ�w�g���G���О��k��Q�Mb�[A��J��nO|���`9T��b�+�'���
UF͋/h����S��V�L/�L�>��ڪ�YX�����;��h���'03���2�2��f��b2gz1�j�T�%��ҥ�\y���e�% �?��Z�cde�듴i���Y��1�>��U��\��EB1�����BnQ�z���k�&F���'m�]q�w����FOU	ޛ��k��'/w2dW!Q,�;��vq|W���|��Z�\^�>���oź����N�� ("M���QEa�v=@�?�0���T��S�!�,��.�赩����Y����� �a�R����g��o�]`H�c ��)z�=7�:�/#ڝ7�7Gz� ���kg�L*!�÷Rw<G�S��lsa�����&#����ޝ�X��[N��,R��]H
&0e��%�X?Id3ũ#ҋ�~���PCt^���2
���Y�҄$���u���(9�"�.�ژ/�P+I)aCPܑ�6��7P��jp߫���e�F(Z~v؟� d^�X�9�iⷄ1���I�H����	��z�i4#/��K�6���ds�)�2�ѭ��\"��岭�N��&XO+#�>���A����O3���tLh���j��hƑ�Ij-�|w�-$b��|�ݻ%�\��ٶH4�(mH�U�0��H�]9S���k��.���a���X��]�3?_U��XE��D��v���A%�D�ۦX$  �N�j��R�� d��B,d)��n���Ѡ"�R�_l��`hG~s��f`ў�j/�$UkrFv�C鯃��t*Rl��8��ڔ�gD�Օ�	aK���M���Af�FEɴ�b��ĻSh(��A�6����K�)8d��O��A&1
����-����T���"zF�o%���΍39T�����uF�pt�a�ȇ����[!-f!���E����VDι��F��!n&bC�%�:�q�7���{UJXB��?>������� �Ӣ��2����
�B��T�G�RE`���h�^ 4!X�_��w��a�k ��Z]Pb٥��������n�\]ס�hʊ��n*\��K1�0 ����12.?�J�?�xHy�^h�|[& �Xo\�j;K�_>0we�ǯD���go7g��lm���\�+�7�;��9:r��E:1���vJ uF��,k���刷�FCJ�������'ZYZgoގ/�K�O/�ܟD�`�V�~G3$H�3'^�V)B?��7�N����՝�z� ��A�ihk�����Aݼl����$e��]7���7'(ڲ1�������e�E(�+0u�%�J~�cPj��ᘉp��+��a�(����d�����\D� �����l˘0��a��-e�V'���Q�������"�M�b~蟑ϡ|��dm��|�2�l�(hq��?$ ��S�[����b�p�\f�gLa��s���* �O_�t������<���>��K���P�={{��q��<aoA���^�3i �X�:v93��!Tz��=-(@JS�H�!k|�ʫ�!{�w��e�֮�A�41��+��0bxG�m"����m"H����"�z"[&��VL��z�!�άܝ系(�!$����}�7 �Zo��Qvk����F�r� ?���>��KL����&���9��Qn)$�-������[�X1�]�I�-L�TwT���_y�ߚ#�iT�V�{H�}�1�r[G4��X���aC��ǉ6��|!�n�3.Ǎ4E��rd�%`��9�P��s8���aK*��&�lؠ�MV���\�I���"ִ��+�2�_�xJ���,"�W)��'HW����o���GrCv�spP�Sl�����p1Η��6��$�%L5�ux�����8���+F�$e��"m���W#�G���{.Q
 ��T��s6�r���$#��z��2o�5j�Z���X�i*aD4cr�#��O�X�2"r�k·����`���2�J�y�l���o�9H+1oИ9���Ka%���hm�� u�%~2�lS�ڼG�l�ulf�G�9g!���R�����ɪq�l,����C4��J;�u]����1�^<��/�=tްf�-�YUP�֋[�<J{�Ȗ���O7��F�xŨ&%�oĖE�g��9���p�0�ܤ�$5�����ԺՀ����D�2"�	f�循���y �]��������#R}��k��ߘSjMr�����{�Z:R9`������~��Y�� ���T�̢��d5xb����X�w�m���2����۪�������S�'�X]���7wtNß������m8K۔�-;mg�̤�����:L8� y�G�g��pGU� �73�WV=�Pu��]���%���S�q0��80Z�wF2�bY{T�vL��/�5~O�J�(���<���>G�2)Os��x��m�*�J,�\��Re&�d��-�-����S؟uc�".u4' �+�qWZ��6��7je��{7��[�^:�͞��`�Fƚ;c)��Z�Vʋ�FS,�)ҳ�ݧ��N*F}��{�}�/�M���ͷ
Z��%^H�~!�����d�Y�[�V�XE���ZN��Q6<�i��i��Y/�XY��A��e�w�y�i*��*}��P�]��
��1�r��� ��^ǺS���y�"κ��K��Ž�@z�5ʏ�m�{��eӊ¦���(���g�D��y����Ոٜ`�[������c���/�Q꧳�	(՝*�ԈE�I9�O/�n�7Uu��������3+nl��6��9Z�aF���9��qi�Xc@!| ��I�Q�&��Gp$Y1��a��� ڼᅶ�B��5ٵrQb���C�0��ڥ����2��֔�)1���l�),Ҹz8v���AI����8�K�`	{kg+5�^O��?g/��b^��d�e�!�8�
��Ŋd����q`�lX���������=��N��'�oi߅���^8eVK	������B�x���M��WG+�N����6�����7��Jn���جA��@���Eh0�X/�NϨ�4���b��u��XS�� �D��E�r�_�L���?{�d^[���w5�;������E����-ut���{���(��g���g�{�*o"��2��8vH�G�)���ǏC��s��[33����l'O�<���I�,�.(��&����T/5���0b��'P��K�x�_�.6��C�Ү�Wy�U�ՐFt�H��/�����Xz��͆���^gX`�:�1�+Qo:L"1��x���U��$���Ź�	����_���YpŢ&T���xѽL��,~��-��� �V�5�����py[�h�	_0��|�シ���2n�r������\'���������iFÞ��E�3�g�$K�V��w�X}�>|�6-sc���:��̔|�@XYD�XI�9k�࠸���?����J3z��	 dRdV4Y�pKH�n{i������O�ǎ���!��h0  �t� ���cHV)�%E��{��jMI��ϴ�8�����j-2B�:��]���BgG�&^�ǈ| �Y��}\e�qIF��H(a�z�*���I�����N��4���.��?m(����/����
\l>>ZcPHE�犪O���!0m�{�dq�Ji�,�X������G�O�uT1�q��Z���`��)
,u����������m�~���l~�}�!d7�>uv��Ɵ��Ku�)B�	��99n�0���M��c�8i�d'	��z��w�I���,��ц`x"�1�����ǣ�B>�����:s�6�E2������{G�ю�A#��f��{�b��P:5g�����M��$��E���b 4��e��B4��q���RA��G�zG��F-��x ���Ȫ�$)W������3\�/QA���9R��&�a���a��4�yd��!�+%?�m��=�_'�/A]�7%��'/8��#'U�ڌ7

�E�|��u�!_3`܎�t�da�\DqCd��9��u܁���*�s����Gu.�gě�GB�G�e�4fl�kv��@̜�Rȏ��5���L4�>���f��>nI����>�E�e��+�u��c_?R�0y����ɤW������:��RlȘ�[��O(�H/r�\��^�D�,HK�(�׈0�~ɹϾ�p����+�����]E^���W��|c;^l��<8��TTGv=$��uB/ r��gL7��>��k���%fΧhÅQ'(߱@��$Š~�ّJ�a��j�}�*?�5h�&X@؋3�s��0e@���N+O���>��$�?�S�� �4��GA7+¢LIHBu^$�$#ײ�_Yk��+W�%{�[{���	�n3(���!m�E�oH��R3���O��O�JÌ�B�s�*���f�7d�%��d��(���p��R꒤�;�~W �J����*��Q�h�B&���u\�+��$��[o\���g�ȮP�M���4e}&��u��@�Ia/�7�
$��&˟�Q�v�̰����bt͙\�xK��N��}��nR��(1b_��V/b�y�� ��n��m4��h�7�7N�w^���r���Hu�%ʤ3�hԆ9�����6��1�W�Eh�m��^��)"ތ~�_ś��~�
lq< ���T�H���2�$`Bgq��qL#e�3D��0x�J�zZ��-�ސ��Lc�RKWp�.��{�J$�*~ݨ�I��B̉�a'�O��7� �Z�.�^z~�U�OI?�%��{d��S7S����w�^�ho�^q�@��/��-�;&j�vZ�/�mÔ�9�ˑ��{��b����>ja�;��(��y?�י`��%Uyz۬g��7�6�H��9�@/��cDB��g�-��ݲ;�����0.�|����d���'� G��/��b�� S�Sj��WK�N"%9V�ys���QIw0b���fW躔M��`bQ�&w���|�\�Wj���a=a��ډ�[�R����|��Q$���ȣ�cGXDm����V/{��İ��[���Ε��*=`���+��9����|Q+ҥ��-?���b4�E}����.� �Ѩ���_�ԁ窇��Kӡ ��y�%�p�ULxL3��Q?�T�[�TҶ��1Z(���H7���;��M�Ghz���HY��e��Iq��N*�ȹ��K�����J�3 ���&�۞ŗb�1 5u��({m�T�뎬>�@��rR4:9�౦���h{���g���T�`�+=.j�D��1$�G[�4��V�Sɗ��ռ:��	�t�+ڟ-�W*ըX��w�]���mc��6<����recQ���

��Y@�Lߠ��;F�Y}�,\J�C R�֒�YS,�v8Q���ڷ�x)ύ3IY���#?M�Ɛ�m扄-oO �9n�3��I.������AiJF�>��߁|������)���j/�m�5c���i���i/6��h����t���,:'�b�-HZ~�^��8��s����0�`��6�5��v��#q�:�l����֩��PHG���5#ℴ���h�'Ɏ��bF�U����&�qJ�ىv�%Uin9h�q�{���1���w{�L�_h_�݌B��p�w=�k(r?j}T�V����pbPh~� ��݅��#���(.1f��$ܸ��򤪎��Hra~=��׺$�3��W(I�O:?.z��ܯs�c������[�r:�%��퉸l��D.�6*8e~tYӆe�[H7m���>�X�?5��uO)9΂��|2�R�W�{NȌ��Rf>�Q�W/��ds�FzZ��0���)���e�W�b+�v>���IA黈6�x�y�ۘ�������}��� �m�i���O *g�(p��I��o��_	g��Σr1���Kۛ�eX����;�,N�e������H��t�����"���X���Ȍ7�)׸Ð��X��9�^q�:�Ze	Eλ�_�wx87����+��BGGݽH��2]D9|�3)s�iO*�i6���X��J�}�{��	d �UM���4�'�I����uU���K�s5G()�Ve�0byط~G������?�ϐ;�"ؖw؜ㅛ�	��e6�g�IU&.�&v�qj�k�� �C�%Jj��k����ζ��af�o[@SJ�k��H�Z�s\�*�;����z�#�+��h�w��<�D��$ p�z�w�Qv��	��VWp�d��e5w#j�)���謆C��*o@��T�⥬p@Ӫ}�%*�<�CSs��\ɒx���ܐo!����uYgq��1�p���c4��^O�}}V���<_�k�>3F%-���&�9�� � 	H,����].���܂���Z&� v7����9����7_��, ��XYd�
�^�Hmک0�gbfn��0d�O�ڱN�ZP,\�	�1�b���M�4K-f��B"Z��&)�
g����H!���}�	�t%�Hآ�+lQ�C�:{�ͻ��Vk����,aI6�}~����]by�mhy�����*��U�Xv���<p���J�BNʠvl�#�g���s�)��`�)�������~88Ty��m�Ҽ��IMVU�I8�VI��(�)�(��w� �_���%/ߏ"��o� 0?nz��tN�o���)�/+o�&P�)̽/�X���d�u�����5����!���A%�]9�O��:!��
�p����<aE�M�_��k�@�au�z��orn��Jz�
t�
b9�a��D]���M��ini�8eX;��eѷ0?!u�\؝�Ƃ�V�g�+�Zy~ET շ����pxz���Ԩ�38�,d����Hf!x��ˢ��	���)�b���0�sE��.���K(�F&\�оrH��[ioJYc2~O�2o������3����m��v8��ig\��:L /����p՜�DB�_���7�V��"��*�4櫧�M{YI��j�L,�h+F��}�_���yg�`,}K}m����؅�^Z$%��Ҹ�om���b�9����w�nJB/μu�Fp�>�h��[w� �78��-�2���}��a�s��=�N��`���%-����0ë3��|��-Y#M�l���S�C%}�A�����J�����]��Zq%X�;��S��T� �n�"ך�jMo��k�x7�_f��������!\��%�`V+]�S�V�7����a@�;h��k>��q��0����I�V�e���&D6Ц�U!8|��K�U�1���̗O�{�i�� �m�#hFY���:���x���[�!%���nZ�%6�� �Q���u��1�`�@������`�\c^& K>:@R<HH�!A�t3QV��_|��}�P�SMQ5�j���`-L�̤�b��6RAĳ�p]S8�����`��"�a���>�vvrfRu|^z�2����UD��+�6�ɬ��U֡�� "��z�ɝ�U�����E}�{�M���}�YU��#㉟@H(�J�U9��ܤ7"Ɂ2�B�\��o����Y�ٻJ��/���޿ⷸ�V������#�Q��sfQ��^$��1k���I0��%�yK�d>�����*����d�N��/�FvB�\��\�'1B����TYS�N9�]�|l���P�?]�)^GZ�E�
��BȂ���|�~o��S�v��acT���#���mL-!�L�E*�*����R���c�.Y��������!�̎��Co0�t�!���xv� ����jBQ��a|v�L��?��ͫ<�x��(�����z�Qkj��n���P��|#,����\�x��~L�y�t�����r� �c.߻��B���s�0�#���º�q�R�͢���� d<��_�o*��H�J�i���1ͬ�s�X��>� c��мa@��Y5��g�bd�Cg����'&P�]��I�^��7԰W���PGXS�p�ː�`��4��z����n/���(�7�&8G�sӢ���f���Z0A����C
п!�(M1��&���3���	z��x��R��C�'�ߤw'#�PU՝���iʙ~����A��mw�~�:�2�{i��C�Bޫ�z���%��� �j��W��`~�Ѝ��Ϧ��03���pn|�٦��;5mY|�>P�*�%P٥b�s�Y��h���P�6�vR��wȉ8T�F{��v�������JIR'?��P�XPMT��-��"��MҜONU����5��z*����&�jۅc�ee�`�V�x��cz�7��K�� ��n���j&%&�� n������&���n�	�<#�5����ܟ���Rf~a�zKQ,����/wW@�A:���q�&��P7-�M����m��{ �vHtL}2̀KX�qu߯<���o��d��Zڲ��H�f��?��E� ��}Ϸo\_M�:�P@)֫����_�DS��aɋ�]X%��Ӎ^�B�����K�<rns�[ߴ�g��I���`de�Ƞ�6�{�����Y�Oқ�����ΪFd��wJ�!��=X�7&զ�c��R��~��.�ٴ�}�q�vꢱ�R��3k)�uCݩ��g��-�{�j�����)r�R	����*��cV�E����zauwĒn�a���9��
Ӭ�4��~�G)F��%A�AI��=��cJ��U=� k�j_s�Wb��D�-T��H�̚�RB t���_h������o�����x��Ձ�L?x߀�	r!��%��m�%2��Vi�y��H�(��P�)��[���J4�6�p��C�N܍u ٝ��& ��KM�u	z"ړi��K�n�Z��=h��������O�:%69����ְ	8�	�j?X���G}���X�H<�x��z�[�T�S��.���?��y?��B$@X�7��=�=�Q���9��f��"��7'u�wNd~)j`����gH�~T�&�-�ד�։�Ke��U�g����xp3i00
7/���9�/7<�%��Y
����v�I���]8p��Qo�L+�|���'��7�0sZ���
��ST��˫Y7l�]�6�F#�.���O@��EK�b@��m�W^7w	��Qݐ^/v����f� ~��vs@.̖��	D�˻@�Bi �J1k�k�|��M�'Ԉa
14zjc�M j���$��PÊ�p�DZ׬Z�U����-��2���'��J�P��N���d�'��8�,�K�u�qƬ�:Au��j�R���w�D��:[uW�ț+�������}/�PFZ.��σ�	�f�T�rQ g��ӑ�E�`@�~��,_���ge[K��Mf�r]5���aǱE��e��8�l�	�<�p9�I�E�K��(��7���ĺ9ʈ�C|����!�l�Л	.�1���h�#������o�`�9�$}�^�I�@gP!��X��mjY^$�N�2���_2�<-��7ܒ� ����>�!G�Q��s�v8�߻��{�Sv%��b�v2���a���
��|�k�x+�`���!�!8��ǅ��v{%c�m����(���+�؉,iՑ��� 43s�l�kJ����ݼ�ą �h\�!ǶMZk�|��{u��3��8aVE�;V84��L����:ӗU��*ӧ&����Na���-��cU����ɥ�|�U߃/	T����t�h���1Z>�g�>��wn�J�QݟL6s��$�'T;�b�� *3I3�4<���0��\n��\h ����F�է��Ջi����4�`�~���y��3�qnI\�Y���6�����K>_�|*�,D��D�Xp&�T2L� =J����{�Z�0�idQ��E&���=i��H蹣��B�B��4hs��]�L,Q��[���[F.�ҋ��M�賩Jm b1X��� qT�)�H���Nq\���������9���QŃ���d��&+�!�� ��t"9��+<@h�W`mڕ�}/ULA<���3v��k�	宄<K�ׂ�XQ ��K��G���M.m�'�k?r-e�{�[褲�=�S!ESOӇ�3`������DMj��'��e���.�-گ�y�M��|8+^���	�?��iD���ن�5Lo�WKBXLr$�~�HNHxiɔg��t4��N��������
o����䪽��{�eMLu���A�yu[⟘�4d[K�����׼44�_�t�Ω�I4��K<�r����P�X��C^�Vz��[T��ʵ�eWn�߅JG�9K:Jas� e��)Tn��n�������)��%����2/���8W^�k�����ݝ�M�CEG�B��Z��|�� �!�66��whs/]̎Js ��Z(js�ɁR�,�pc'�;��s�o�:�ذ�M�v?���C����.�.�Κس'w�U�"h/6T�b�_�폓����t�W!�8�I�\��8�fѤƲ����(�X�~�NÔ��N��oۓ2��\�ۋֿ�IQN����<U_DFV���9�ӈo29�~_[|3�-z�e��l��L�{��}FV�9���N��sm�����x��Q��,=Ǒ���� �6�PsR���Lu��$�r��Fŧ_�N�Exd����m*9.w�k`�L�O�� 0�1�l�'q̓��/������� ����!]<H�5��ި�I��^Z���ħ�T�:��,�o�LC4Ni��Dj�x��^Mx��@��&��L�~T��#�!`���0�c�խ&Qv8S��B���G�!ѝM��ϼcnX�� �h�-�_H�p{�\j�$=�˵.���T�.gD�c9��>'Q�I�ȅA[����Oaa�I�����Sգ&�b ����Y����{��[D�C.�IE��������!�b�������Lv��`q!��^?���cS$��� AyL	b�TaU���׉�u����U�(6}���d��߮L��!	8_C�[����b��Q1���P4�t�^�YŁJ� )Cp��I*�� �$�V�����T��+��E<��'0ހ�f2������R���j��[?N�kp���~����d~6vj5�R9�Z�뛳ˎ`!=a�cu���(�q\��k�$o��t����^������ݜi�ș�qƘ�l=Va˖�W8p�)k3S=c�R���I��{]�q��W��U��K�;��J�L[�\HڠJd��t&Ҁ�T�ަd�	�i7zG��bc�3(�c�1�Ҽ�կe��"���G;Z��Go@[�t0e�v�����h�A�td�L��*=�]��01���B�0q)�@��&�$������� Hm_FM�j�.Y��GW���ʵ�#}�@ʳ7��UJ�z�\Qq(�]�{�x��̣v�F���;��y��$x���ڰ�Xi����M�H�y��9� 	�P���.�����m�!�A�^󅄾�٠$�05_i;�.��P�w_�*������ ��k�{?RQ�>���� ��Gp����طhىG�O�\������'��U�-�wSOf/=6�pޅek��������	X���hf��~  �"F��5*E(M��I�l<(kۅ�|-������X���1TT$7�KBtF:F�J�'�ۇ�y9�<��!ː��~T�;1�^��Ͻ��q��RS4A�r��a�t��K��^:�
�HzTBN*�Oé4O�m�U7tP�p ��xUe��LM3g�J���c;�=�}W�)���i�΍D��p����#�W���a����(����`1{�w���VX��A>�|`Ub���*)�Y�f1w�5,�����q��s�,(�[~4�=��]F����19&�Ӿq"�A�&0f�GeE�&u�<�w�J9wcv��]|3���c��$#y�dF�V�Ǥ�s�E��e�:|�^��/�b��-�s� G��I�X�|��Q�wl�,�t�����[��M쳟ܵ��� Z�]���틂�0Z�JT`]��2 wfp���9m���]��q;���!�E��c��ǗQ�F|w�ʖ�o���
�|0<��^V_�����"42ֲ�VG�DE:	���a����5�p�����3�i1_~ ��F��p0<·(��:����&
�j���͞y��{���Y Ls�%��
N�XU���#iG0��fȔ[,��tٰ#�$��J�;깴Z�2���u��-~��E�S�d�D-5�[�&���:YjS�=u_o+�hdd�j��:^�h?�nue��Q3���kob��g��=Mɫ0V�T��nT�����]Ӄd���2i��b�{��[�J�ޱ���}m��p�� �~=� V�&���B����d��n�2"����D�ʐ�:w!56����BƸ�"F\3G���37R�E����� ��\�Q�̩��C��>Â��и	ȓ-��c0�ꚺ��c�2R�je[+���}�4S�E@0E���غ���E�c�ۂ�E)����J�?���n�������k	�����p���4|	�CY���ܺ��)$�t�νh�zڻq/������ʂ��m��Dr�nBRq�����Z|�m���F�%6��Q��Xt��G�d�%�7�땙�+�����d�`z
���(���>��Ny���`+B��1r}��6���A�iZ���r ���Ư���[��,�0��0�sAa��3��#�6b饃R|TF&6OG�>�h	�C9�w�lF��ɱ���HZwC{q+�3�?���C�YmQb���X�E{#$,��+�0"��{M��24�wP�,tj�|5]B}�X�� n�H�b�e�uА�g%��$���,*c۷	J���� �{��n����K�aOx�<#B�%ʇ�Oτp��f(t��Ĳ��U9*Y7^.L�<eX�n����P�syx�3�U��bne���[���c����ϫ�ғ�]��g�� 6L�wM������o� {�����揧���c�댏g���L)��5�(�U�]k�z��e���ډ��Ed����)0[1W�^�c��A���K12R��8%oP"{/��+vX��yo��-R`gY�T�^���/��L����,�9AJP�q:���p���7G�q:���>P/�D,���:��)V���zh�,i���$.4t×����\����8���w�8��}�Y�Nצ����~qؒ �.i#-%p����1�A�8E�2܊�Ŷ+o���ׇ	�ς[��.�Y&K�Ko��\OG������3���i��p{��o�=	q��`V#a�w���@ɺ��P�p����Ö�v��m��D�B"� {�5���\Tdd�W$�8VJDy=�xBn�������[)�r.]2j���k���O�n��㸹7a��BNu|nQ�Vv�H�<.6khaX�F����H���28dJ,T��ؔ�5���G5�҆���;�h�M�Ik���5*]��Ӭ��qmG[{��861yњϧ�\�y�����u72O�����y/�*e6�_q���o�=66��1R�v�iQ���/�ԑf�eS�J�ev�*�efDp:�����i��?[y�!$�K7��ʼȌ��t�b4��d�;g��X4�@̓�Eon���GR��"5�5�!�����- �gz.��`����I���~C�-K8��)�MƊ@|>d.�-)X6>q��Ȝ��l'����o�!�P���#�H���/�)�ͨ���M�pD~��1����v�Y��]5�&�j�tA&Tk>��̑�8RhI�(\r(� f����N���E\2�פ����	���M��ժi��*��
���&"ˍ����a��_�ɾ�O��Yơ�����q����\�탐OO�T�t(3 �"�#�TUR#�v'�;uc�f��$�o��.����B4-����h
��*,�U+�x�Z�عh�U�GMrb�+GyA�wƴt���"�f3+��v�2�`I���zߥ���w�O�I�z�H�;�y�چ�,{��J͓R���y%�!�ۓ=�|	��ap�׮ �"�m^�.��d"S^"
S�B�M�����h|�e){�0��ʗ��X�n̄'�Tn��[��A�m�[g���|YfF�ҦO�'���M�{�	��궙�b�)����G~�+EJ�]T;�;4�PN�]�ws6����: ��}�w�m�dq�|9��\Hŝ&�\s��%���W_��]ѐU��N�)]R'��~3���f��cڋ��n�83� �4�xY| ���*�w~��ߏݍ�C��9
\vtY[�������7|��hw��$�FgBo-UKpj7rt�I3/9��pj�p�z��g��lm�4�m�HZJ����wD��=jmp�sO���i�>��f���Z�D���Dn��ף6<��')�,��*큔�o�:�֤�ƅ!Q�^��2
����#m�6vpi�s-f�ӮΘQ�k�����@3�+���#-�tU��@��?i�V#V
��Z�CF~�u(+�V����VʍC��.��I,�k/����� zK�N[����L:�׵��m�xi����zi�>.�:�T��ZT����<`�(�Z�.ҭeq
·B�b�,Dꁭ��u�`�x���ވW����
��e |��+vs3G�5��[�3��J��������@Wc+vpM�� '�j7,���*�m�؎����2��W���^5��?^�<U����w׳i�����J8J{>3\��3+�֐��ު�zJ�~�
�z��c��B���C������_�.�x=;ّo�B�(��S���?�YE�]@�k�/��e�2�f�{<&�}���v�K�V��y�a@{�x���/��Ar�so���S���Խ���*�W�,�3�ܞ�������W1�C?*��U U6^)(��p��;����P�uw%]s￺�󚰜!�=�6��~<��T����ޠ�\On�M���^�A�	I	�~��(m��l*FP�^��e�3���L9�]�
i�����n�K��ka�Ҥ�P��i�d�wso%�<�t�wE�c�39?��U���e�{�x�g����β���-_�@�¨�$�p��G9���=I�$�~%�2G��P�aY�[!cG�0Yv����Qz=;�
����
M��8eKY��o��[�����>�Lq��cb����(qhJ��p���>����=�[����/[�:="UC7�7{�a��@h	!���^�[{��=��h��(HD��`$t�=<՚�ʍ���YNӕ$�z*��{���#}&S�3����H���E�U���nR-�_��7��L�{�^�_�����wn�hA>ku��~W�����,#f�S��u'A�U��+ �9���5Lp�|���H�~DĜM���l���h[�@t��V��*n��l����d���'@wNè*��f41�',O; ����}��B309[���q,���r$�"��/�UM�q�t�j�t���q�$(u��'��an��.XW6d�zޘ�j��;��_u�QH�Ev�_u��ib�@�d�~�L����^l������m���<d�Ofz/�$�9�Y?���x(B'~��e��v:ŮY��z��C|�N�m"a_�mlD/��7]�p���L�d�:p�[ύ���3�K�O"=R8��<����/�ف�.���;z�!�~m�_	�ܯraP��i6j9
jr�@��q-{�~hc�_<�ƨ+<�ɧ> 5/�ZΪʜւ� ����N�.њ��O�ՠ��s������w�4���mKt-�rG@�{%��%��\�+3Qn;^6�!���2۠{`n �$x���g�����y��e���"Z�'���#X�� ��C��p���̪`EL��?��I����w#!�b0J�{U�$5{WT���X	�E�@x9�G,���Ƞ�̈���TCIk��o��
����$��?�t��/�E_���O_�3�Zȵ����VPL����~��1�� /�t�������X�{�;#!+�I�r��0�n�IbS����".�dﳌ!�a��D[rW�m
+����i�p��9�1�KJV� �~��Z�R�u+�{��Xn��`-�j��eRfy\T��x���akN�>�+5S`��5��q�lg��.zs����k� @J�}���XF#רo��ݟڦs�M�����ᦐm���Qp����ɘ9�NP�+`տ��֬���Z;RE&�������B��0?|A����6Ϩ�tF<�#k��5����N����R�f�T���)A�޼.��`��&���D�S w�1�p�"�j�[�@\m:��.l�H����Q���`?&���Mκre�ԣ~P��Z��Ӆc�e�ލd�O�nM���q*����§Y^���d>��Sv�(�\"�\��|���@0���-\�yS�^�+g;�8���(�P홀�T����S�ۇ���Ǫ��\AVT����a��@�#�U�D?�[�S!��򸴭/;�	���|���'a�鮯~cC~���u�b��?��?�ڬ�n!��������F�~('��&Jv&ib���F���,��zح�7��K�E����W#2�-s��|,�`H<'�vD�g]���,nTlSt|���vs��ޏ�F�u��7��դ�r��i-���I�@ �u'%}w���(��z"rg�:(�u�cn#m)n���;���F7u٫��6�t��>
7���L>�J�Y�fhql��2U��%ż>xv����~h��a��L�����9C���H��v��;��\(>��28ȪԦ����tm@q����)}F�Z{�;��z~�����a�hp�/�v����-��7�m�B����&�&��[dY�ǁ��b�F�6�,D���Z�ר��ߛ�'��'5�R���]�3��������[��[���O�,]�pۤ��8��,�i��s�/:&���8��y�*��Q�aC��"I>֖��j[������O�V	�|W�@`���,�N���5�t"b"K0^��q��Ia�~K��q��nk���S���.ۇE��Ҹa=����]#������9z2m��x�X]jH�j����u�����h �!d��;ք�)8Dg���r��)��9��sEȊXB�W���mfy���,�ټ�KF�*��5�}G��D],f �i��^��Ժ��O#R���4ٻ=���i��� �_�3@g�qU
�:"���w��Lh�!h�u�:vb���:�����]ë�lF��Յ��X�,y4�[dpf)�@qCL6["2ґ续��6��9��i=^a�`�l�8T۹���q$2���ݒb�zo6	B�����B�Z������@��$b��)����/�bmK쏺����Χ3@r�`��O�{6�*Rp����%!��K�w#�d#��jA�6��[��U7*��v����5��5���T�a��k����:L��
�O��_,�W.�,��Z�7�r����d>��XH�����	xY�����B^d�l�"@����&�R�IKeXwH�U9���J�ɛs���N���EM����N'd;p��CkiRbu�eP%�31�([nH��k|۶���ɯ������66�����D�oң��`�B������UF\�]���U/�]O���1�k[i���Y ���_�hg��|]���o�����')�7����E�J�̿Q�D⠋��=�?i����X��M�b�V���H�Pr��_#��c]�g�_��vm.{��z7�|_�1.�b�@@�6��,�7'}���jfS�e
���&wgF�53gL�eA�>�>�!
�*�;�F������2>�b���VED)�l�lȕr���(S�EYF��=��K�1%�X��ӎ�f}������э/�%�*�#ci��AX}gr%>k!��K��EC}��o���P}��y~�.��
~�phT��>�� 0��wkȑ�9��Ժj2m�mq	�I����>�PL�Q �D�'���H����D�:0��p�\���4u�x+$iཎa�[���S|��o����BT>=��\h���FK(7�.���b��g�!:��)��yF�)`)`��5	�f���,Rh�6�հ9�~��%�d���c���@�*s8� *���kiv�9�sTg=���㩵���{Z���t�R�����T-&�Ѳ��8�u�⦁lH-�F^j�iG(N������y��,�*Yun���_u�o�H�E�#��Z�c;E��2�b�����T-%9#p0�q��5�0Z�K�J����
��x����an�w�~/;��4d���U���(�kC��?6$�Ù�ͦ�(�܃�eα�Y�]	]ΰ74H`��ï�(VӉ]zq���A��\��>PM��AdZdd��Z�}�Z�*:����h��#��l� ��Y^��k��w�_7n���'&({��_3?cWn�OD�����W�FA�SqŲa}�p��0Ϡ�����9*�0��p��b�/�Ȫ��������_���A�
gގ�Ec���L�F�IXJ��|�,1�XR;���]P.8�YhHo*���:}�g��JZ�g�D�$�Ɲ��#ٽ{B��(�~�`�����֙����F�ݎ����*�W��i�v;��e8<�Ak�}0�N�6G	���<E�6Q��O��٢������"0���	�Szco���s�2SG�����XD#�.+���&���r�	�5�;��t������k4��)��6��r�"�p�A1�yæ��XQ�,M��ٌe��{���)�_�[M%\��{�>�E��G�21]ͮ2k �JD�b�\�E�Zt7�&1��iwU��V���Zy�n� +Z�{[K����2������X��ю�E�ʆ�SL}~��ޒH��{|b���'B�[k� �� �.��VG�k)Irظ*A�a����ɉ����F�F�m�!�W�d!��?HQ��2:�����7M5*�/�� �n�$'m�i1p{6��Y�%�+zJ��N��B!$�*��5����-):�	���UN.V��hO�x�%���gW"�]Y��,i9roR���=�V2 �2���|Qv�F�W�ME�$E�}�(|����:"���b�룮�]�J��@�@� o]#�9e��+A�a2�V��昶Lg�yj����ع\���H��y.ܐZ�Π�I;�9{����RC@Q�nxs��]:���;�$��_P���k*�[��g�U�����d)髌9�Md��Osy?eU��?���g��W�őp�ڍ��od���j`�G.���ϦvAz��$�Q��4yt�֑�$��ψg'�'5�y��w�l�ZC�1����v^X�9���TU��8��O�S�SG|Z��j��YpDfL@� ܈.IS�-�z�'J��M2�"���^^�]o����9k��͐Vr��IPmD��y�1�ӡ�����B�G�-إ ���P�>DX���m��.��p+�V�J�V�>�μ��>n��m�Y�6xh��٥A��S~�ߏ"��PЙ\����G���C:W��~[_vQ�6i���tdD�3�IlpH`�:w.Q�dg&cH%���h���>�����ǳ��k����:������t���(��%)$��h_�⥕�>�b������n�g��|v�Ϙ����4V�,��X~�	z��(�g
me��(W3�캎Q��ޟ�ݾ`��\��\X;���D`�8�^����@�S':����kX�>�p�V:�P�Go�7���s�G�� 0�FX���8������$��B��d�O�V}ޢ����� +��[�"~8.���ᵏ3
��By������E�t���k�]M�]
=��<��;|�\!�l�Мк��;`��]K���k���Q�WfoIS��%V71d���a��^aa��6j;�+���9���M���""�#
��� /im�HD5�R������)">x��dvo\P�K�p��ޘ^U��#���(8��{�KO���x�s,���D��ӇV��D9�e�.�#��1�i�Z��p/�]���=�;�&�5;
]d�Y�t˳C��ۖ�9 �_N�ELn1�����<k���\��>Bg���I�_��bŞw�ގ���}�x���W��W�'���l
�c9x �È�6X�aLT��¦j;qGV����g�2ۦD_��C��y�5�ke��a�S�[vu��p !�/ӫ�@h��|��)a�_��:'T~���w����!�}�e�Ŧ��K�Rmd�DG@ټ�v����E�&�R0Q�:C{m���6#O�Y�^��A�	�4��{��Z_g����k�ޅ�n���K�@FI3t���F�ƣ���Khg��M!��<_�&II���sMі<?���]!o�}S�f��Ō��}��t���
.���$}�0�c|�ut�FܸL��K\�AHd#?�#�ԅ����w�� .aXg1��
Ja�u��r�}��_�>0���ɳ�2'Og��S��a]�xk���}�fu�]��?@�;6�Q���"V�i�ɪ����]Gw$�SʬR�9h#����е�VWd�����;�(��*A@s#���0��IpW�����
�	i�َL]:��5��Jty���˺ �'�+|�1遗́���2+�7����+�F^ހ�le����r�<hh����Y;C��3iՌ�L�D��p�4�^h;���#�m��s����"c��JI�P(���g�ހ� 1|�����Vm�ܹB�0�n����o�2\J�x���f3�\P�S4�у����&;�qo�G�Y� �iQ$�l��tD�c.آV0`��9?J�7X
�۝��e��&�1��z��(vp�����,ӧs����h��J#��t��"���%͒�ʕ��>L4�Y����4�F���/+��WB�7+���㘏�@�,P�y#�&�Q{�Ɖ�>�B�ԾjS��7m.�g��<?2���V�dl7`r�R��}e,>��	h���]��T���2��)U�����ՠ�,WzקuXa��P���)����'m�ڄjٗ�/��lN9,�Я�Qج�c��n*���F����(&��\;�+8ፚڻ��s�@mP1���:(��ھt�m�C����Q����+��L^��"��X(��Fa��Ԫ�_�Uכ׆֑,Z���g��s���P$�]{h5}�X��{��$ܴ����#!Ru���K7J���l��5b� ���w}_��������F)~�[��L�5��pp��Al�l�D!���6m&���*�P�7�!�K���4%7�q�@�%�[��/�.o��q���k�I�S�Uçm�>�j�$���x ծ79�)���uWi��SFY �M�.
���Ga����Z��կ�K�}-/�[�^�7�v��m�j����	���s� �5#�\�$�D76���m�=��:,�M8g.���;���o���_m�ajM��Ó��+X��/>:�sZ�JʨU=���;_/�yp���=�>�������+����ͽ���h���	zHQ�c�Sں��̽���B�T����*��7�M���8�<��-�
9���$�Q��9�U�h��]qEEh�hQD�
5��.�m�<��J3y��)�t��xh4��,��d��A��	�V�(7�es��bܙx�!C��̅gk��0>�8��n��EQ�y󭽳U�n��Q@�]F�w�	�5���κe���/��&��$i���~��N�x�ʇA���\���%���ݝ >���&&/�,Vᒵ�r�(���&P[/��x��XA_xP�҇O��P-����V����r:�UE��e����)��*q��,W	Y!a��IO���(v�՗��\�W�^��"��4_� ��Vھ,c'�Og�h�B*�.������-���z�:����=ݾ�?�f���h�&9���LV����oG����3�g�7Ĕe=���4�OAh�-�'�z�&�𮵵�< D��H�����̓�X_.S��r�l
0�VVɅ�]��@|=��{$���tx�LQ�1��.���k��#���d)�iAC�
<K#S����D|=<7L�B�3�Ax�f�$����U욅�`(�w�uư\8a&V�!r "�A��Q�X�	��j0�(\��霄�I'��6�j�2����c,�.s�\�;c�rl� ���� �CU3Nm���#FV�}b�:�K�(w�XF��2?�1��c鼸��t�N���ssa;h��D�R#A���;�+s��$��)�ƎƆ��;!�m��d1���Qun�H���J	��>��_r�S�|���F�%	��%P ��6(�����fӑ�W,#�~��5(��