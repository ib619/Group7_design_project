��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��o�Y{NĖˬ���P/{��$�)f�Y㈎����� �9H$������,�-_6��6t�y
�ߋ�M��� �����J����)S�r�P%���xn���� �B�!�93�e��$e��X��v}�5b���\[̒S��*e��f�j �S`M�	W����}��b��4����������r(���=
C5���Z
=��������
�#K#)�ʮ��K��%��ƒGb��`x������)�6�5��y���z;ܳk:��/y`�.��,�O�	�m��?�PH���B J����-�f��T���|R��@nU�>��ЦLG'��	���M��N��߇]�.�Y�~�tL�����_���h�W�l���]}�J��.x`"��`kk��T@�t�)J�pߒ<96^ʚ+S���_й�]K�~V3�jF{���a7C|Ĵ�W�S���I�5�Z���:	�c7+�:1x��M�d�[��2�v��=��?��@���Na��ʲ�+��zi{�p��yy��%��G.JR:J't�Q�z?�zN��{���y���=��I[�~�e�4���w�^
�;Jo���gK�9��A��>��+&|�P� G6��a�˓�?��-�ù��+���<.�2b��Ƿ��&�q�d>�_��.���H��gCU�xYPэ� K)��7 3"��Qb���*U]I�B��/P�V
$���3*��9C�N-@�~F��#sH�Sb)���:������hQ	Bo��>pˌ�<'ګ���B��(s �;��jPK��l��XFn�-}��y�|�$����v;=�P��q�o˃[��pv���g�4��CL�H1�4��0^�F
�����t��k|����8�d��*_ �NUU^ٗ�J���;���c͊�9PI$'׈�?{�4�
K2d�ۣ��r���g�a���V��h5؝����@w��k� ڡv�o�
q��)��-Ұ�U�4H] ^�p	�˃���b8hs�o�3�G�-,+���/HY�Gފ�<�򌾎���wC�$C���]�7S(R���������O"�T�8$�3�5R����NQQ2X��78��6�G�t3�K��8ODk/҇��7K�L�ѡ�ȣ�
�o����fH�-<��)�_uNt�ǧx��ǭ,�ab2ݥ���1� �b�H湻�΃PՂ�đ�{�lRj( �5���
[+c}�Z�i6�:r��$9��k`jv�1�?!�;��t�$O��/�Q�t�ﴣM��sd�$�����
^�s� �lM�M�h�4)H,ԗ�t�T��`����Sa�E�41 �(u�<�}��$��,��/&��D���~0��l˖��<P08l
�Z��F�j���J5`Y��ά�*�F}]k�������W;o:�6R�*�&����CD��l��Ѯ ������悽Pv�@����7Z����.�VEC�"������p��aN�w�[,Z��}� i:���Y���E�W^U�q�K%,�|����|�G����u�q|x�XBzbQ��R0�j�K�eUKif��*n�+���V����I6Ps�W
?	LG�e�ڋ��"�k��q�'�f �8��싪�J�;��>�h�17��;`i�L�B���^گeUj�h�Ƈ�Y�s����[���܇m)�Ѓ2��;�zE����"X�w_
��A{�^޸1��-	��/���=pb�.�SO�p��m���l��a��^6�+�Fcu}Wq�a�h���=��b��h��ʸ}�s���{�Y��!4�Zxq+�{.>{����67��?^�_p����m,e��ݰ�L6a������-E]��ޚY�������i��B� m�����Ԯ�c҄���xǉ��N�c�rU}+�aqƦ�>a��;����9}K[##��8�6��j^q~
�~*�Y���R�
��qd�>�< �w�s�c�������t�H0�\�~kr2�>U�\�k�$�ݮRi�f��"Q��5O�SƲ�C񯒸����?'�؋?��Fؕz�cCe��[����f���A�э�u��"����L�M���+#����l��M�Z�#藎 "�jb7���Xt҆J�O��VW�Xf yu�˦��O�k��l�^�I�Y��Z��^@�4���.y��Z�U��l���jCCa_�na�MH�fgv�E�JBP%�Ӌ����0V��z�������L��d|�~A�R*%)��B�b�OD7˅��a+_�:DS��;h_{Y�K�}�gS��α=]�[��}k�屴Ar���j�c�ٷ�$i�scF�qC�bq�kf���.;����.�V����j�R��fW�^���@�� x�|��\�.}��C8>�@��<�x�J�����Gz�lk��+L5�]��t�3:f��5"�`:�f6N��P�yX_2�����}�
/6h?��#�V���r;��a�	����$��dv�;�+U3ML�Ye{�i�1E���Y�42������35SK�f���\��T���Pa��~W������!��D��T�;��.��+ژ���&c��o�S�z��^C��(*u�h4u��;�.� �	��2��a�Џ~6��,����qy��
 ب-E=��Cв�w#x��j��_RD�d�y�iX%H�:ъ!1��g'G0�ߧ�c�P�/"���E�A����{�>��0��Z#���-�
������l�9a�+�W�Y�4�8�)#�MT�՝Ɲ8Y:-�y^�>|��=��3e���ڡ��-0�/7�_R#��ɓ"<�pE�aKS����4&�.i�~��c���r F�;e�c���!�Q�� �H�٫,�0��
�1��M��i"i���jn��!�#�@^�o'ݭ��
�rM���������m�
�m���\�%R��s�r�@BO&�Vfj2[UE]�4R��a��?�]G!�r$v
�2��۔21�N��� /��2\�(�i��� (��:^M��?ն���4�/:-�"�C��VӬ؇�횬U��v
�hΣu�!��ֹU�KW��I�1�u��k�g���Z�fj�|�k0�+���)��܎�h�n�����K�S<�5|�}�ً�#o���������!��^`���``i���E�K��<���ͤ��d0q����?���R�qs�`���/6$�Z�9~����#)�e�8��Nځ�j��/�Tl��X4U�m�3�����(��g��
_6Ѱ���>#�Z�Y�'P��7B0 ō��B {|�:��?�f�k�W�~�@��i_2�=�"}��1M�.o���^$�Oo$-�7�T����?=7PܮN
¯��1��ޜ��9���kI�Cw*זk�r"�	u�BH���M%���j9H��"�� ��Ԕ��ڡe�'��0)��=h���e��ނ����J����皆@n�K
[����H�d?�i5\�G�&�����qb����70|����y��g��L-B���~�*�1,���l�����B�u㝛��W����,5p���z��Ͼ/�@�p�2��h��U�V`��'nԲ�Y�׼P�4��x.[�ڞ��Q��rj����j���3ADC��q�$��������wH�����ս��m� a��w��-[��D�m�q��_�SM'�TJB��He�QV;5L.��Q�c^Cve�	u	�gSN��f�h$�d����96 �!^��"]]s�[��b�ǃ�D�R5Tj��_������C!�1��yEY`��(2�Ա}��-�AFZ�:����R���9���D$ޟ'H��^~q7�^���M�d��c��+k�V::��e��u&b�d���ҥ����V��H���Z�����<L.��*F��bm���1��t�l�YD��%e8��+����mK����h�mz����ՈT�g�y[��$!�%;p���j�s�c��������i����G�A8s%!��Yn] �Q��@J�:��R� ��al���ǽO#zi��I�^/���yu?,�ёB��b�Kl��Qon��Z�ZKD���dgb��A��z�D
�*F��W]r'�[��
�k������h ;*�X�h5��@�1�rC��\Zĭ��%	lѱ���$�?V(�p{'�b��w�{�i�>��Z���`���=�3[%)�<n��QܩQ�O�z�X�ь��j]���~�'X/�3O�C8�R�K~���0 t�Q-�GY��%_D���