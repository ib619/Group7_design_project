��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p�8�&����b�B�
���:w���w'y�GO���w=���Ȫ)K��S��.�5��Qo�.v����I��D'��El����4�@���P�RG�ERC������(��_���Iv�{���E�.wc�����x=a���v-Wv2zo���	��)B��|�P-���ɺC@B�'#iU�Rx�k&��A����T�-����@ه:ɳ�@� (���#����?�ڎ���y@�`t�f�KzV��Q3�@��ʒA�f�ĳ��Gz�uؤ�!��2�j���\�$QF�18��!w�-��0�a�Kr�o$�� r1�(�#�"ov����[�F�Z�O�{T��g�1m$�[�6B�.�H>��@D*�2�޹mFCu׳�B� �Fi�Ƿ.a�x�H�u��ƱM�0��Q��%���z�83�����:�ɾYϷ�4���i?��'����2�._�$BM�3�Q������L���� c �2����SԐ���r{���0Z���x�v�0Y�C�JB����)p�ے��e�ԲlH��<��
V��̚�r緥�IF��DI��B�>�7�U*C]��3B2H¼oz�S`n?��$Z���q�K�c`��?�3>�����}=O6��x���צ�7i�s��8������7�����N�.tS'"ň8�$J�)�t�W�B\�����Q��{��:�v���n�.G��&��I��x/���u�z�ˎ�u�n��bx/a�=槅��$N�lp������^�T1�������}�������0�!E
��7��7��R<G�,dEyWKd��l��*r;m�������~�<SDq�,eG~?���l�<��PƔ����������j��CM�aߡRse�fu#��93��2D�.�%�/���V5��	�nR��;��K_����o?�1M�J����-oL��/BU��p���5Kp]�[H�����X`�B���ZCJ*�9���xH��!�l���Ԩ��>��w%jS묞\D�4�k�U�=�؆D�2^حɺ��t1�6�����v���h
)�qlm��?6��}ocR�]͈ۋ�ں#Uw�S���ɋ�!7+Ƚ�P4aaZ1��,u)�l!z��lq��.,�ם�)#����"=���*�t��*�Z�e|�$f�#�.���NY�ō����R���ź��/[������v
k��4E�	��b.\� ˥��7c�T�bP����Xl�KZ�ҫAnF_EKEy�X!�}�Է?�G
�)T���w�6�Z=�\�f���#��U��`�4�G^b��F��B�[g����/�J�l�� ����c�'�b�U�Ϯѡ��!L���.�_z�KYTKTMM ��8u��߫+=o}vb��adY[)��=[�	��>�@��z��0��4M��c�0,�*�Iڻ�S�n$���B�K(d�&���ZA�1��m�xa�_�'�I��R#c��߁��/�����j �X�I��=����9~�� cRjI�fO:�2�>�^�v�B��3c�L��Fȶo�X8�Tc�t@��:��^r �Ж'Q� �2"U��œF���*��`��pB�˼��"vx&b�AG7�t�0�?����3���> ڋ��7�*gg �8��1"~��G(]��7Eȃ�ꯏ,V�<�pi���0e��p;yq�щa�\u:~⺿LL�3h�o������dQ�.D�ҥ% �[u�����m��o5z�h�+�ߊm��j����O�/A+�����k!q�1��"�%��)$��g�$ �;8Z{M�BݦK��c��.�8r���Ň��2(�M���)!�ooϦD�6�U�~tSܓʙg�ٙbv���Ł(��3�[n3���>��u*��
�Mf�/�J`b���'^��d���L�xL5�L��iԨ��Ո��A7m����e�)wsNv�yRo�~go�0&���$�I"�� -'f�(�xv�e��= ���҆�'%qx�<�d��{�ζ����43��`�/�I�u�p��"0g�S�Rwex���c�ˉ��vO��UCxx]�}�R-��d��&%y�>�ȱy���6�b`!���ެ�]��pa��3�z��	L����x޽h��z�)!X��P��h��z}�S�6���tW���/��ɝ�V̨O�~D�[�"�>m��e0����P�λ�:��e���C ��Lpv!W��6�-ԟaq���J�~��&����?k���A��>�厛~�o��(�g=��*T߄^c����F���>��%Ei�Q� �)-\�˞ߥx���x�q�j����/cI��>���+1�����^����;�%O���=o��ȍ۳��߯�"��eW������+���3/�����j�*��R�Wȯ��W6���i�ۿ�q��~�=�}W��Ȉu�������c1#��~f�U����Oɔ,d�*��J�y�MD<6[�z��K7�ev���K�o獁M��1"4�H�?1pkpk�N��T��.�bަ���S�M��J�H�|���������Xzt�(��6��թ=gQĪ�����<r�����޾9��G�9��o݈��Oh�p}#�E)���Wr��/�nv��|]�H��]1�lON�-�r��T�����"O�%^��B��	liv�ys�C��6E�MW4Xz�a�l�^b�p"�N�O��R��K֐��5��'~�`^%�׳v�j�*b���"�'�x�}�1}���0HN�.C�d�A�9�] y�**5C�C	��h%S�9�Kd��AuHmyă<RÀ�8b��#[�K4����w+옉�3*$���fV!�Wdބ�0�ͧ���<����>;�v~��f�pwS(h0=�l7ٽ�3	���`9�Ld�W0Z��n��}ruAo(�ů��_���,����SAҷ��%F�O���H���	�P�m�[.�{�ӕ��⠥\�D�=2�/��~fH�b�_`��s2�U�3�̜~�P�%�JG���cI��,v�i�Q��,In�.�ƚ��ɢ��9��>(R�V?s!�`1�|I�m8����%��>��#��-R=�!7�,��>��#��j���{d��5ɾ8�?���O猀���z1@�a�WG�ШCA�/��N�Jb��/�O��:'�>э�F�]�\�)K��"�Ltr�ƭ���5GN���CЏ
�xL5�!��;��eMUK��%�@�\?ܙ�7DNH�d�d��D�V�!���:[H�0��b����(w��N�y�TgOiZ2Y_iV]��߲�iu��B��1�,���+��*,g�-��~���S�+u)j����G�5�:*V����E�/U�����`T���z��Lq��T#B��5�c=G<�5e�Ks���������c��B_E+��H|�Qo�v�v dy�uI�"�LnRꠖ)D	5��^h�Ǭڔq`�L���� d��T��87�z����D������i��?L�j�]ㆹ_8��y�bI%�M�Mh��`��%��I!'���06ٸ�86��$��=�NmQH��O Ջ���(�*Υ�q�P����	]Dͯ�T�(HK�񂘈��(�W�BV2um�`:��qDa>�I��p�9;e*s���||��EC��("���"�'-�)�#��`U2G�ڑ^~�'#�����	R�!���m��B�u8�sE`\/٤r�΢�`^"��nP{�3�d�FY'0`�*/,U��ɒ� �pl����l�k[k����'�c�;��p��f�����>4�b$�@;�g�&�ŕ�}�l�����>z������o�"���.��c�̧��|�Gp�?��"� H�{k-�R��x�!X@�'�a�Jjp��Aq>����XWg�6T:���G�����ڒ�&it��i}r�3�X}͐��u�:M'k�]SQϊ���X �������B,@����<�����I�JK��oq��|��*���t��|��H-�t�tN����6w���S��_vL1e�M�tS��*_U[������jt��~�h΋v�ChVd�3s���D:��'�t@e5[�An���x���+���A~_g�ê7QQ��I�`�C5Pw�W�8�<��d�H4��frX!.�Y@� ��_���Ʒ��Y����UB2!��g��$�b��0�W��-ߙ�����~���)����wsLB��*�L�X�2-o�Kߖ�E�t	����� 
�s�ǧ��+WS٦��P�ق�.7�Lwp��vĐ�3]�e����Zc~ct!:��Ć��ʰ�y{�/�F����ʮd�=�Ĥe0@�2t,e]_	F����R�/��r�_1�V�l�T�O��/�1�XW�)`��m��W
I�w�ӫQ��P-1Iܻ0<�$��Fq3�׹ù���;@l1ճ�`��g$��>��~�4Vű�u�����9n�|t�0$�@̝2���7��ֳ�y��?�^�)g�z�G�N�V�J�����P��J��?�w%l�`�o�3 ]f�����s�\=��-N�"�L���в-,�|��nM]�H��t	���s4��)'d�9#}�L̎ ���6I~sI���]��q�fUn&V�#҂^(�O��@���6;�sy�>�aa�쎻��*'ΈQ ��Q*�\54o8�$��'���I�i�Խ���fmk�k�WwIĸ..9Q0P�[�A�6ԈX�%H����S�G��&FSq��7�%� ��Ep�f�D��Ƚ6��$!G%�8�R8tl�o$-u\���76��D��ᩦ@X��|ڋ��&�W�a�<���&�΁ǣ	O˾޷�.@�O�8q�xd�;JnQr����VKx���R8��x wr7��)LyR�oĵz�>���o�*B7D�#[X�(e1m/=��ema(�/ ��"�ַ�P>�ֳ	ɑ�o��&GO��G�+na/F�y6p������0Ƶ�?Zb󻕛�@�9��U�����^~�U�-���}�$��Vf�K=��|�E����3��>>O��#����=�+�¿����xﶼ@�S��*�W�,�Ж��xF� ��~�;�X���u*ˈKL�7���f�9ݗf(��Z62|�H៱^��w;䔝1v�{ш�'lX���8��+�2;������W4Y�{.	�Y�+��$�ZF$�ôF��%�ӏT)����Kb��&���.�u��[���Pf�l�ӹS��7�2 ��t�����m�A�)��)Zԇ�߀E��Ί�;ซ�dsAҧ��0��`?��"z���=g��?�BÓD��}��وR�L=��O���3���EP7��IϽ��7
��\KA��~��n5���?�ب$�9A
���k�K�8�$��8@&oW�2����ܗ9�� ��_8�$D��G襃"��(�i����T�φ���m��C��|�
uC��{��x{�m[f ��۸A��(��U�i��]֌a�t:�37aB=��BzF8ƔOe��Q����H��o�\��i��2���������!��{�$�pF┌�͊��ё��5�K�h�GB8��3��U�e����VI�G�K�>�}�U��C}�eqqFj����d�u��B��o����~��Z��+�h�Hp"��0�����}# �DLa��c<��l����
�mO�F����G����BZ6m����԰1jq�)���*DG��@��4?2�7L�g�;`���3�L�X��ѭ��ܜ��W�d�}"Jת�M�,��t��r�I���$��Q_V��r�,s1koQh2��',� � x���l^4�Ӭ@�/�`&O�y�LE��_�w*�F�T��'�R�b��taA0�^��F� .�I�Qc*��������v �}��<�i�[�*F�!���"�C��4\Ӳ���]�� R�]�t�_T������;ku��t�͒0E���`x<��Y�GKc�Ȉk�!�C"7���d5 �v�5��S�O_Qi�3��"
��/>w�
n�]D��9�P�O��dp���憖M��>2��m��d��E�BX�i0��r<�X�8 ��(m*}$�F.��MB�No�%���?��7^ ���!�eU�1�s�������ؚu���SE̳_�
P�%?�]0�\0��%�����i_�iP4ʡ��t�L�k(K�X�!�\�o��)H��>�"����K�H�D�p�d(z8O�gN�|��|s�Z�2Y�7������xZ0j�ee��O���@��٨D��u$�v�B�ÛOTc�?�Mba�!�]�_��D�ֆ�Nrc�ϱ�N ���*я���E�\�4�_l�`݄�C�$�E��h�3���c&R�,�U@4l��刨`�BB���У�"�}�0bL�
���f<>��v�>|)ܬt�n獌0��^��W��`�8�W�z�8�'@Q0|W��ޭ��K/ZA���<?Z60�x˓7��Zs?c��6E���L��-����#��[�5$����.�C��1@S'�K?-[��Xa*�n�}~�<�3|���,:��x��+�e��N4�*O���:d���C�<cc��G�d�& �U�U�l��`^Y��{/3غ����[�ң�]�R��+�'�i�ϗ���P��bvI����h��oO,��~4���`Pތ~b�$�w�x6k�6�##(�m�����G��{F���f8�+O�9ׂ�4+(`W�@��(�st�0���O��e�Nb�'�%_�0��,�M�Kw5l��jxk�fJs��j|r���]#�`΂�&�:2���n�)�������|���Sc��x�樛�@P�:�.΂�9�?Hy���Y����qP4h;?��:�S��u�j�>:�����Z�p$Ko?�[?z�d���m���fX+sbw� �=\��O��G4@Ne�@k�E�jqU��w��s����-@Ֆ�zK4��H�7Ei��!ujķ�?�;D�簽�8q�h��e��H�P5�p��'��-�{̊��_2`�<���n���������$!����%7�eX_\Y8��`6R"���2O'�̭�0{���en��6�}�����0��~�h^"ۿU�R����Ⱥ�E�w���r���)v�^*唪��z���CiEo�N�˷���%tW ۡ���dO&Ea��FOՇ"j���j���#U�Ō��܂���E�Z߳}�w-W�랳��
��R1�LM��.Q�P㈦���f&)[m��<UP�c�K�=�z�Y����P�Ӫ��Y�V���4�9y���n|u����0bn�YM�{	��?�;���~r�&y��ꀯ�CdT���2���!��f��r�A:��(��tC�����F��&n�iĒ+ն�"ai�_e�&�YT���5~��2�3JQ�s��;���fe���kr=�8B��S��