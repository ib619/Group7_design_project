��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+p��F悢��o�Y{NĖˬ���P/{��$�)f�Y㈎����� �9H$������,�-_6IX$�������ˬ�Zn��B�k��b�H)7b�WˠUe��Ǵ��A�VP0�0��{ߤ\z�ύᙉF˘y؍�����
����;����k�j��F����H��ja
�P��QK�悅��5�sʮ*q^���lF&��OG_�l�ic:ɽ�.9x��}=f��,aFz�:w�;��E��L����^q�j�k��5RBl���XN �\���a�Tr��kR�5�A��yQ�^f�n�ȇ�I)���;��~�xM!�ԧ=$�z�c����s~@�n߳1�����顭��*Ȃ�!����Ӑ�,��D��
z�@R���ڨ�0`|�Р�ڂZ��y���Տ���K�9� g��ėABĎw���"�� p�c��r9cqGdsA1R32���D�f	��Ț*��j��֔����w%s0?��O��!w1��ȴ���4��0�K����*wϒ��r��@|wH����@G�����}of�N�|�1j��!��q���O��oP�@���Z£v�u���?���<�󦏌�C���p�9C�N.���Y���?��&^��yg���emɵyC
Ծ�E��S3�[)���"�߰�;Wąι����)e�A�'��p��z͕vv�Z�'�~���
v�;�2F��MA�h�x3���Fצ9ਕ.�7��@"�����Ӱw�H�7�)�.�ш�/,��h�n������s����*Ǿ��di���՜5�W~�D��I�;Ĺ���\2�]�j���8#k���:�o:fL�ج��n-���J��DC���J�6Ш���Y>��A�蜲::��yK�T{��|�ۛ�/���-��F�Wއrz��3u��ɯ�/㧇�����K�#�Q"ش�j�& ����K�`�é��QV����l�(]���-�K��-d�S��O������Lӵ>������ݘ>`��Rhx���Bt��序A<:�ߘ���Q\?쑩� ����ݚ�#�ơ	���8/[nDએ�@H��CI?F�F}����_C.�6�s�~*��]��U+ ��j���X�={��v7~�AE!�΅S�T.��
{U�RfxWzjTT�'��o�M�.g�.\���F�x�>�� 0�tn.�"+��q\ڹ�9��4¸Y��Dt����R} }͏�Y�6e?ڴ=��*&��f��VwVgz��d����g����h��M�߳�3���\c�~C]��
�9<��O�u-r�i�M��j�>ɀ4[{X�����MD	��|"Η���l�H,�bsǜ�O��Q*,>Ū�Y�HUt�W�����/Ꜩ�@p�U F��v���jJrho+�h槳w�T��Ɲx�^�l�	SW)���=���b�#���f��
����xQq��z�� ��[�	$��k ];s&�O����F~S����*��wp�$#����C0����sƪd;;�7�u?r �C7�Kۂ�2���-�r�-�Ns�Ǧ�h ��d�N��e��®,o#p_�]��aq��ϋ˸�n�IL�|�.�$�J$�I��:fbV\5�cu��Ve�O��zK:��kp,}.j;0�_��`Q��+x=xd:�\`L�(Zg!�ढ़pR���?��!�L�k,�B�
�7�������j*���M�P�����<����L����~)@�|��7�dg<p��g�02Ǝ«�s�\4�2�y�� 7��}3�9u}`C�}�ߟ��9RH����K,4D�(=4�']r���1�g��h2�y�s�+�D������/�ߘ�jb_�͢��qg��#S�ǰ |�������������0��5^tD��w37�Cبk�(��k���1njKb�wZq�,p �6�ye,��Q��`p,v��l��^�g��~wL����U|�c;�iI�''w������2:N�tK���&g�I�P�x7�+�P�j�ʂٛ-2ǫ��'��Z[���a���TA+��ܨĺۂ"��nds�b���Q���(`�A�.1���L
�!�V?�g���R!t�9�[u�p��펼�y�n88_^��e;K�i��U�y��1i�r��#qx��ĭP�pߺb��%����zت5&.�d�(걃�F^B��'�͘4�����a�q�&��3�!<ÑG�?f�+Ќd��jO�g{f�	��$�������׏��1�#`���0�o��oI�P1B���i�*��1�m�k�4���AO�2a�9�W�*C���՞ߧ�Q3l���<�?>���3�zK�W{L�%SG���>�"^]�6��\��&ě����ܶKf�����&&؁:m�e�.t@u味k�?��z�+ݱ$���B��*��.U.r�󾘼+��8���)eט��*W��F5�N82Vߞҥh{/�	n[�@��)�q�~%�@V���A��&i�v�e����*!�Oz�ΙRP$�ͼ9b���$Q��bN�#*z�u� 	�}%��#�hザ��
�mݭ�.�5ʬN31s��0ᦇ�Ha*J�N:��~҉��X݈w?H���1�n�B��	m����(�Ťݑ�$K���̈́�؞�����t9�*m� Q�{�C8���;�ocw��9��2h�5���>M1�xs���'o4�1�«��T��S�"g��:��>Ar���!АMa�Қ���!���G�Ǹ���y��\�0��q��~d�3g|`�9����~dY׈�@��Ѷ�^��A`���es��
�a>��4�#F�4k��b��Ѿ���䋔߆|rd[xs{��Y$���	�I�
�U<S����f�j��S`���z�	�� �z��	a�HL?�+SD2�a����t�Zo
B�����'�]W֦d>��tU�\��z��r����/:D~2��2L
*�'��Y�0�q�,h��XSw盾o�_B�@�B&���$z��D*:'�P/�~�;�!K/GI
�� �|X0��X��!������Q�x�j�����ግ54���y����loѓĳ�M%��-%��y�(<B��T$��#:�t�NMJV��,sͅ���:�jW���d.�u�՜v���m'�+Eh�D����؟J���O�#���1�%�%��QS�ؔ���~U2oH�M~Y"�*d���QG����U�S��#e��B���j5�#��r`����ƎNoе٣����b�[=g���ܔ��V��"�G�˔{rG���5��V}�i�⊡� �fJ�k�'���qv����<B��;N`�� �?bh3��y�=^y���*%K�zD�Z1{���{��h}�\2IR!��ZUk�D���͆���HU��sA{=�J)1�z*���<�}}i�%�s��G{����gף�,|6V>]��������t���u����_��Sn��f�'B��JŃEj�M��
�g����� �o��!�(grʃ"L�l��e�M�B�>㶈j�%)�LM�yl�C�Z�#0���8�dz���W9��`~*����_q
��G�ɾ��,Z�y�ay	���͗�*�� ��1���&�,hZ���$	�J̧D`���1m�$&���]��b���@=D�"�C�#��`ٳ���i�v���j�\L�#}D���M|�a��#���V7c_!9=�,e��s�(l��dOh��O��;�0WE@�D����$˱Y���o�!��k+1���E���'� �@���x��� ݛ�\;V���gYly֩D�U;��h((�[T��K5�^�KP���9��uZ���D&,�"���`i�5��b�T�%S�T,��zz�]X�d��Y�u��s�dm'Q!7[(eŦ�htR=���BY����;?�!��I��Zy:0��/�4�����k-49~ק��|d'�2�_�y$��ș������i�������=�+7#L���q��N}Q�!�	�+*̑���^D:�%h$�l�d_��ɝj�7>�˿�{%���x�fi��C��8%�z���W\g��_�/�y����NN}�ӳ2w��*6���o6gz�7�|��×�$�
>Q��@��k���Z\W��2��Ѥ�������j��>��K8-�H�(�߱
�@ ����"�x_���V�ک�7&��]m���4{iT?ұ#P?# ���K� vՃ���l4��K��Pn(�|z�ė�����>A
�ɷƪ�ػ���.��������p�*�J�+��l,�9�{����iY�c�sw�'�Rkf�Ɋ���.�l@~���N�i/�1��C�m��`W��]K̀�j�Ù�n�����K+=:2X���A� ���'���aF$�7@���4[��|�ϙ�0h_�^�Dwv��-��P@�AU�3���(��{,3�]�? �E�ȑ*og��K-���w��*�|p��$��5�:wed���Ȭ�<��`�����-��!�F�"BF���bq�e��R�t�^.\�#	e��&��F�Wh�޸�2�,��sH�"���lQ��dI.q\���w��{��i%k�L�xq���q���^3���Fp��
�?�~�}��Ԭ$Qr	親��D���S��T<��ϰ�b%=�bb���&{_(O��,W9~%~�f���<�w�H�� qTJ�H�E)/�"��X��K�y��E�zF��k�t��ĝb����\�=a����#mzi��5���^��5�G���u�{�U]�w��x���q����`����J���2��
��yNp^*#Gq��䳗#��#��mzM�&TSU�������Vo�>.��L`�S�3_�E��Q5�z��2�<�jVT�` �Oe�%p�ug%�j:�'VQ�*3�����z��þ���pdɇ
0��	v�����f���E뺾�U̮u�Ų6�oY���-�EQ�qfF+GN�	r�k�6#��a�d�x�V���smG����؁؀�������c�)�>W������3�B&�ٷ?eZ��7���t�.j��(H�����$���%V�F��}�~%y��$���.z����ڣ/W���d5�݊�#��r ����rS���n>�lF�)��ߦ���z��e�T�}p���FCim���3]����Ȩ9	y���F��M��",��-4�G[D��r|
B�5t�,jJ)�,��HQ��b������(�g�R$�H7�8�`����Į�Xq�̊Ќ���/�r��b�qbv|���a�R�,\Y�g�@�ͣ�,��l"���.�L�q{���l��M��H�����ꦁ��`�'x+?�w�w��6ϵ�x��kb�b���~��6���fZa��K��N��DA�1�O������޷G8J���nGx�=Ҳ�'���J��%���
�z�>s��GD�޹�6@a���^0���`6F;QG�a���>��)C����n�r*�H	�>��{��ϒ��	�o7~�ɘ�USZ��q��ѱ��~O��|�H��ʣ�����.��Fv�3k�J�hB�.���4_��$�Aƙ�[���Xp.ߑ��Y�P���#m�'0����Y��C��<\�DOd�č�o�O�"�N�}n�O,�^��r�\����{r�qg!xe`�]��QM��Gx�Jn3p@��p.�J�|CS�e� �z���:�8a�9:��_H[�Y�4fn3�f��s*���x}~x]G���Y��n�&�c���x��$��'�8hs���S�P���x���I�af�3�E����ՏȖKtpm�Aׁ5�*E|OQ��ګ&�ˮ��,�r)%DG�Ǘ)��l�(��23S����F��K�0T���fž5�B��e��a:��6�ͫ�,�aI*��V
YQ�o�.��ד��B�������ԜeQb�AA��E������!�ɶ+f���AB�/��x���I����%�g�d��+$�����BDD
�֩���7(]R¡��@3�L@]��O1_�]���b��L�Ŀ���[mَP�c@k�@d�U6��Mn�N�n�^�h*��ؑ?���4����u�:�c�̰+O��P]��U�tW*� ��Fcɵ���,;�G.�{��$�Nx��_.#8�-'3�?R�S��U6]� ��B��eb���'�".�	U��I� ?f�8��Q�,����AľðP��Lr�-��zb:	VV���m) ��mY߈O�pB�pfE�\ Ol�G)T�B�d-ހ侟!����Fzk�w��e��q�.̿f36��Ro�������<S�0`��6F��kј4�g�N;o�L���b%��P_��>�:"��?�dqz6>�*�&
h�	KP��M��t�ѸR{��pO�x�h�+÷������/Bw��7���fv�MƱ��U��e_�H߫��_�o2��}�6�i�bJ8���!���=h�A1�<{Ot�w�,��)��]���Қ�B���ka���WO�����;u��՟����2#,��Z����XN�Ԫ�BE�͸kSp��h�� ��(M� ᭢�֍[	I���@��fvژd_���e���\-H�ulw�L�5:����0H_����ENJ;�s�B΃P}FFB���c*�u��g�!g��Z��-�Gc�@�Ѵ���)���8q�n���[V�!��	�s]P8��v����1��fV����{<jլ�[�3��R�4ܿ�����2������QV��&���T�;��P�2&�s��a�.~u<���CC���u���>\4��-'	��GcY:+���a<�~^�d�q_k��"V0z΍�1��-��b� f���s��>±pÐ��y��[Ōw,�z�pP��xSeMOr���[�-Y.j�G�vO�^�cu��:��	��ܸ��]�o���Y2��ׁ��iՂ���w���8�@"?�(�I�~�h���O9B�� �'�� Z�,s�/:v1�~�{6Tk2OJ� !ك�o�rLε�L@=�X��wX��7 T۝�mO���E�U�"�"�9v+.��)�kROC��u��6g`��,ԃ�tKFӠ���1�Ha�L����RF�����@�ه�Zm��9��'��*�t:N?W���{�؋^~�U^r�h��=N�����(/W&��e�U�Gu���ݚQ��(_������� �VCL�t�}� tk2y�Z|�09��pr0�R9[�S��p��A�>^�ڷ�?��VF<,�0�kls�.cizu>��<�jG�V�3S]t �,&�=��Z哓v/�6����c�;�l��}�vg���"6'A�ǜR����7	Nn�N>.2^�W����n���:�D��8�*�K�W���Q�@Y���]p{�9�+�!�FV�qQ)����ϴ�Z��gp� 	�y�3\RU��ha��%�,RD�s��iB���Wa��QQl^��P�tX ?�� .�:�S�p�x���S�@�H��j��!
�l�'�@�}I��7�e�*"�.�s۔��gD��N��xܒC��dq٨���Su֐Ʈ���ݞ�zr:Sq}����[�i�}џ/�FV�Q��f�|�O��Q�fe�S�UR��2�m�grĔ2�߰�'������
�4��sC{-�z��메��M��>�[N����vg�2���^]��S�7���k§p�zP;�����'�q��L�e�K�oB� pu�V��E��YV'PL�r
n̢���c�E�9�4�i�UO}��}�aV���W�Pcv9���r���0����#n2��R6>�0��?�~���~gJ��b'Н��~X$��ɤE1K�1�
p slw}acN%
��'�0�#�TS�,�X�C:�u�H��Ƒ�uT�Y�5r�F,�!��(�c�^�x(�F�5��5*a�!7�y�� �P]��C]EĹM�W�����Eѭ0�f��l�R�H���j�Nv����M����ds�/-����)���|D�<Xx*���@�I�����ن}p!�����nv�eӚ�yP��b��=
�a�|HO�D _qN��j�s@m����Sp
K�8R��ŵ�Q�B�Ft������7�-�@T�B���ҥPtV�^�~� ѢU��S%�{�F`�)���K���UZ�NCgK=�`����G����ا����>��#S&7��
��{�J�\��!l|E
3�Z�k���l�B������I)��0��<q����`L�g��D�L�� �Q ���tиu+Ֆ�PBiU&��qN����tL�[0�kc�IATW�F����)�D�=�
�E^�P�ha%�!��o���M��j�%І��w/A�ac�6~ּ����%���#Eo�>f;l`|0O��v�������(UgO6|��*�i�A���R����&���z.��v���t���-k�5z�'�7)"���S�%JR��X����*�R�=t{��Bu
�� ��_�4����Itr(i�#�K��B�]wc������H,��]��_�'O�*��;wbl*k?�?�/�Ge����l���@�uU�@q��D�x�Aa]��G��` ���b�'�I���ҹI�oS&�""mp,���9D_�\��򛧌{0"�H�����f�����/�+D��T.p��Wt�e1H
����q�;��x���sc����\Fu�н_Al,	.o��^H�%t��"�$Y7p^����z|�t/(j��׵E])s�LӠw��J�����]m}�<�{�r*���gH�Ҝ 4v����1�w���V��i���`�����8�N�aZ,Fj�&%��OZ�k��ՋB'$ߘ9���p|:;![�����^��9�޹ǥ�:�1֫ثT(q���ahr|�h��3+v�_ީ��X��4��`���;U3�3SN$�wy#/q�{�9l��g,�A�I	T���K ����9Λ�3�m���J�b�5����������Y����[j
T���B���꣼RY`M�M"� ���@�`(%[Ag�0������`۱��n��m�8�\�PX̑~S�JuT\I�(�e�p[vM}��Q���/��ߟn*|0ߩ2����8{x�Z���R �yA��ÔR���V(k�~��i�&l�y�Ql3>m�)�Te�Y�{����W�O�������Kz?��q��#>�|E��L��*��M�{G����h���k�g��T�DE>\@U�Ә�7�'Œ��Hi]�KeQг��k����,�W�U�Vm�����'�'�Rչ�����[1�󿂍w���\p;��)����X[Π�P�ø@�2���>�j� �Z@�Lq/�G#d,@��Ni�ע
�][F_��iFJ��jFs#5|�O�8k�ym���3�&ia+&I	����2f�v��o��Yp�8��G��+�F�|[�9���0��|�����x F~6)� <��fx��K.��ʨ<����2�A�Q�$�/���9�늗Ԥ���yj��B���(TC��ljR._�*���)�a?�Fg�@�^Lo�]��D�l������v,�#ϒ�f�H߽�-��yU�}*��M8�>��
�'0	��2 ��Q:Wb�^��F_+1���q+�����,��'�J�^{�&� t�PD,? �8!]����XQ*���eS&yL�5Q<�Fb���#+d*.d��[���U\u3��i&-�k���&�n�,_Ɂ��d�~�:�����5�7N0o��n����Ϫ�������U	���|�W�;�ND뀸�酂�H���ڿ�K0��^y���HP����z^�X����˘�V$*/�x�Y��,�I����Q��Z&/99�aGFΈU�05��o��s�O�D������.�$���#3�̮V`ڮ��愋�)ɳ��k*0��n,�]S?w�%��|&gr:�x#�MM(,t^ڀA��Ӱy���q��ؠK�l����d�	�w���x͒�������}��'G&�������T3���&�6'+����ب'�Z�Q����̮:@X���FP���F�� �Az�;��4�Nv��|�0#�~�b�kR�"l�yM>������f#C2q�)�q��q�i�Qfe����4#�H(�.��(k|�+2kt3�����ܐ�4'0�W/K�:<B��{�߶�0�u��4��I�T��('w��n��#q �/ޜ׷�|�x���W�'?���Y&Hp��bW!q���I4AađaȘ�h��O<��+���B�Ƶ�0:LG$�V䅮j2L�P�7W��7mid;d�c���9M�j�l�GH"�\��}b�޻
�eB�+�C�N_(@��o@âb��Tr�=R��7)Tv�	���*Z�?�1u������~!��`�s��7���R虣�5����a���?\�����(&u�πz@W<�.ڗ�뤽�<i�~;:��՝�E7A������26�9��6V�݋�k� ��]hB�ɜs��E���slY�7�~7Ժ�.���gK,,�Ƃ�m9@*"6�.�O��e��py��yg��D��B^�:鍈�az^��/���%AU<Q������+�W	qH���.&��c���m���d�[\pu3���6��T{�2�e)��_��Hy�f��og�%蕍���;6�|�� ;�� |�pI��c�Q�$ی��iƁڼm�<b�B�ʜ���`����~�����b�pδ��6�s�}C�O_�t"\&�a��R	�*�سqһ���Tuj�T�_("���J+��5T^����ǈ���>�=/��A��~u�~[E��T�$R�=wH9oOl�(B�˗��V�Vr�K�o�*NŦ���l�F_��0�fF��\�d���`�5ZQ���٤?�7l�پH�dʑ��ޘ��|�O
���m	�X���5��<� ��K-=A:Kɳ��N �NX�]�.	�}|8���b�.P�B����D�*���b_e��y��� �����tB��"#��O��H���B�	M�FXVE�ƛ�+эL��ˢUkI~���h�o�*?}k�ɻ�"� ֋� �'��^S>	�M�8�e��#(��e��
Ixll�~���3ّ����3pWHW{<p�q�������v�u���;�g��R�_��e�� ��S�Zϐ.B�OGjX0"��&-��7��X�DwF!�"�U���{T�˪,�
���v���z]�>%������v0��1*����y.�W��+H�_����yz��핀��O��@�&��n@����q�f�w&Vx�6���:ch�[���2�3WG��>�:7#��E���z�ݠ��W�w�>[2���,�9�V��jA�J����>hs[�L/@E
�1u��hq��L)�Ņ�;Ϩ亠��͒�AF�0����\�gs\��D�6;�������/2�_�Šlu9��[Yד����i���e(��-����Z�)e[��vP�T��x+��lAU�q�u��k�ov�u�[��D ����-b�N�'�\`�cǷ��Ro4�����+�X�	���f���ѧ�/�P=��j�Y�#�$V�����	<꽆��Or��
C,�ĞC���]���N�y�4,x�.4�c�i�"s��x��1��5��("hN��/Jf�a�[��4��KW\�}���!{�*��`�x�ՓFx �AwƎ�%��"�[.��*ݱp��Ecg��0~���Z�4g3]2��}�Pz�'z��f�Y�N��������?���Qi$��\�tױ�M ۩�+�e�n��P�7C?��|�ػ����{��~ᕼ�.5D����˂�tI�[�8]8�,�_J��M��F��(E���`Z[^Q����{[5@�"O�Ȏ��fN�s�?)ۇ�#9�^�ES�G�}���}Õ���Z��@��ju�aF�Up�Jh
���@���[��y?\�V�\�h0�9w2h���º�٫j��(S��5V^�!/ɼ����'��Z��^N���;-��%#3�4�6o��,b�-��`��T��-M��|�;��}��#���[Z@7�s<"�wQ� 5�&�3'�GS����Z�QV!.2�ʭ�KF^Sc2o�@MQ�zf��9DO�f{(���t74n��,}FqF�OfZ�_aG��Y>GH=$hb��_�������>l������]U��2��Ӊr�]�#��B����i8�܍T �֭��V�-���.��x!��:<t$�"��Ƞ6��������K�����N��e]P4 ϓ�V(��`�ł�I��j8Ōe�������	nKiy!=F˘���'�W8�z ^�x�0'�ǩ:t�Ht�a��3q�|��cs�"/TN{��glπ�
%�9"@����Wq1�mh�����q��a�)&q֥�Au�O����#���/J���qT_����w����Z3@��$Z�P���m���ȸ�*���Gε��2�2E��>@x��i��}_���	