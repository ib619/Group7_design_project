��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��t�x�}�Eg6�3)��I_T���@���B��A�u~1�c�(lW�7ó�I��o(���ت�n�2���ñ���o�!N�Z"���ƛjz��IƟC%?�X��IN]�C9�cYf�o�K�{���V5�h��߽fY_��~HvB|��R���XLl�U�U�Ɠ�iN�[6��&RT��j��"���˧���A��۾��c�����_!�Y�ʊv����;�aԼo��E�,��3��*�V2��� ��A�F��ӽ�P�	�@�#�c��Qܺυ�7���S�J�n�\lBɣ����}��ܶ �9�6��%�Xm����Vq�61l��p����k�X_��yHs���L�iL^R+)��kg�[RE�U�=Ib��xj5~Wt�ufM�L�Gq�֠ͯ���8�^������(�޴]�=��N�s�~�C����E�-Mb��:w1-��;G��m܅���2���W�s��*�R�t��+�!"�^�{iCoN�ȇ�n�䘷HD���#"�]R��G7�� ՈaS�Ur?	�T5�Uwn^����i|޴�`�1�U찿:\�;�p��v��	������hD1ڸ��v�2:�"�e���;�n�[,.'!2����baFԕgM��� S�2��+�\>[�G�kq���L�?b903M��DST?½��}E0&;�F'`�G?ׯ>�W�����o��!��2u'�Ѐ�ccD2ZVm�O�,�}��4���s�u��V��\�`sF��b��g�K�?�>�k�Az�%j=ü1A�$�{!����	 @Fi��	$#�����n��ڣ��"�P圸Ry�����6��߉�sRϥ�-�W=���6�)Q�d��(������[ }�ͷKk@+���ێ���K%ՈP�s��Sؿ���E��7.��9H��F\���0�F H3�y�5���t!�{�vM �l)im������`���X���a�t¦��6'���ƷÊF��݁J�N-�ۮ&��+O���1� �m��4�z㿘�t�vWM�7h�āJ���H�|K��[Y��T��$����)����x�bC��" �N�W��m��^8?n�k�r�`�������n#O����:C2+���k�I͠J��ÆG���56)�g���H�Tc�u;�j�Haw		�	;r��b�%sx]�B�P<�h7}@b�Wv�:���2��5��M���é_:�ș��!Ņf��u����2�	 %��(�(��:D+U+���P\1�,�`z)�rE��B��G� 36oV_�^�ʜ�6e7]��z�5�ncr�e��KqM4�Ь��QBa�8o{��0�s(j��H@�K=��g蒣�%��8��*fYO�u�8�ɢdy�Y��1�)?L���6���qA����G����aֿ�7C�S��ă���N��l��fn���
����O���\$�<�
������Oy&���I>8�n�p$��CX� v�Ej��nq �U]L�.X�K���]��]�ʐO����Hsu"_f�%j�&��.X1��D������T�<��%��ʜ�f�P��9҆p�\Bg�W����ݹS�Q-9��Q���`�Ԟ�؝���<���E���	���E>+]Ö'��\��tx��z�)-]��	����B��%"�C���{'k`�9����'���ſ_g��=�bM������ռeJ��� ��^���ŶX�Pt�{����=�F,c�����_�	v(ю�� �ڱ�O�ޠ��_�yR���جF�1}`_�2W\G � 4�Jbo�ԋ�2oE��O�f�>�;O����U�6�n_!�\ [΀�?�Z��2.]N����iC�1&�7��6v�W���Sqs�=֟�̨P|
@��t�	�%���l�P�����$�!b�f�R���$�Ul�k!�&_��w:n�",u�M�M%E���i;
�ǖ�u#�Hl�b7�u�) ���"�g��); �Ṱzt� ��Z�������	�(��ϞA�9~���uÀ�/L�H�茔�B<�f$�~�`gk�g��L�o��J f����2��C������G�'�K�dDtZ�/h����wT��.Э��<���x��c�sg�	�Wv�H@N\搨/|~���s���1j0�h����W|��*�v@t��&��u<��Tp�¾E����w���p�4�S=�@!dMxe�Or٭68��� AQzh�\�h��k�$7�^�Spm�=�A��i�V���Ϗ 0�d2_���I�$��}�WˮrNܻ�:7���-�k�a�����MR�!�啙1Qb�I����8U��)An��ܟ��[�`6-M)�MУ��Ɉ��S�4e���	qQ�$����YQ(��:��O�Z�F�[{MX	������A��g!�!�C�a���\�bb��8�-�̱�S��(>�%| ��34�iQ��Ct���;�}��ˬ$en��Qs�a�S�`��3Y�i���0\U�׊^_Q>]W�or[Ϗq��ӡ�6Ԉ�J����#��m�+V������p��b.6ܸ}�#��4̏��!V If/�hY:��6�$�<�PJ�;9@���X�{�"p����2jy�O{����D��:W��>\�NN#��N�)���=�EY�lԦ�C�t+8l�iCjy�#7oN�E}U����o�E=[�U���{.��!�Un�n�g|L#RU����66��X�
���� P�G�&�vN'W
�����]��P̾8薝�֌麯�R�Q�^�B��)5"})�@�f��m���y��%��(~?�����y��d�a�	=�w��B�繢�N���
i[�o߆�V��yz�?Ѩ��k�3A*�׀!&�'���F�V�*�-����k��H�0$q�bB&_���) �����x7EhI�4�I5��iF�{`^"�F6�Z���{b�(v��u�m�G�)[Z����gEJ�逡љ� �	�$�,�S[Z���0���hyC�5�_d6�I�I��S��.�'h��<�qR+��YM;�{�W�R�<��5��˗���L�Tr*4����F%�����U��7<�l}-Y������n\ *��m^l�����hƔ���~%_7zǾiY��&�g��iH`pO��g��2�� ���H��WzN ��#�����,�q���&�[k!��r��4AjzR|��.hmpʯ��TK
Qogu�1�4��+k8���P��<"��o��=|\}��71��P&����U�Nh9�͎�,h��vAu�p�B��w�a��b�kL����S;��xw�>����p;c�;�1�F���K��OC�2�y5'W�Rv�nܡ��:���F�O���ϮX)v3Ή�![����f]���Q����|h�i�=!o��@[�6v��GQ;����_C��܅Z��y~��X���ttIP��w�u�ܵ��(n�1÷�@b,\g���A�s9�3�\�� �i䷎�Z׏~���?V	w������Ue��gT�KA���Z��'G�Gdwy�O�>�o�����#�U;�����-�H/ϧ�rJ 6	ed����b�����rL��%���)?�'\�ED`�ov[
Ǒ��-v�w�w$�l�5(�/��%�i��^�P1 c6����6IP�$+>��)��{�����7)������E&�4EnɏR�R��SCBk�b�ﺄ3�iy�;�p�����o�g������*X�B�A_��S���E|wd��gW�w4ݰ�(��/�T|�ԡ#,m2���/��^�z���\��������JJ0�N�w�Kb���4A����f��rp�/���^�Q0�E�����
l����'��&��	6�9�4̚���;Pe�
�m�=�^y�Re?^/-���3T*����������ZDm^����ExK^������	��H�ܐw��g�B禶�W����!	� Q_$}eOX�_��i��n@QV���Av�*�\���E�=m�i���+�%y�|�u�>4^-��|�:��F�%��x���&���M=,�~��\��Nu��25�F�\}� |	.������h���r�;B��`�y��������<a�R��٣Y��Ebb߈(����=��쉫t���s�)~ߕ�A���^k�T����#��Yu�0l:-��\d���%_#�:/��.b��%��]�x��ߏmC,L1��\�����ӌ6�_�[[��y"yGE�5�4�|{qvg�S̜�1���?	쁃�swBi����n������܌a�	�t�n��m����>�GuE��ˊi�ܖ���h�AY�r�<�D%�r�ǆ��Xo�̢l�J)4nx����
< b�K�E���G�?�(�!�n]�)g����j�6�
��U�-�~xC�ZC !b�� ����9�&R��3�}��k2=
W������L�ߧ$�ިب*�:���{�usOb��YUq�`*!�2����p�K���=WY����w������:�\i����4eM�\�z��z	��Ī�?�'"�Dϥ��i�w|["�0�%p�����~R�e���cn�����C�>��G�ދ�w��_d`p�K�n��39��S��Rx�	�b�g�?�e��孉�����5�@�!��3�#�[^1�BѴ�B���y�iɼv�V��F߾	�8�:/ȣ���.?��V��58to2�x|�M��B�6�K���o/1ԵKhD�*�S�%���c���k����hv�������He�'F���A5_f����ǹdh��5����*JI$;QŹK.��Ja���tS�k���N����y]�7)���C����i��-"38�B6�Z�w����)������¦&���E⎂\�Y�H����Rϝ��/��6�XS�����u���
w�0���܃���s�-�tLY%dL��#�T7��
�0���[,��	�8����pVWg]���<��~�/��<	N�(~?�k	����K4c/[�.'o��MD��Y�����إ甌ųfw�����T*�]��/$�"[�6aś�A�7lT7�\@!�H�H4PqM�(��t�������h�7��������~��dڸŷŚ9����u��#��խO�+��f��\Ġs�y���r���r(=X_��%���\���B��M�(��=�)9�܊j-w�e!��d�d�̘�z���N8�~ԕ�W��PF��*:x��kjW} @Pz�i�e^w-Er��U#���'�L� b�T2bEP\G�>ڧ?SD� {!���eT�I9,h�F�yޟt$2q��vi��9���O5;W���:jÓ�	VP���'���Pa 4C�
�]�F1q߿�=~�3z��i��0t�B���H�����$���t7I��,���u������c�e�β�d�I3��Db��d�1��yD+����<�����,N<�u�vC��{.p%�yt��V����\C'v�g����.���Υ˫�@:KP��Q��7��SX*��Ho�Qɼ��p������R>�gyd�����)H#B!{����S��X+(|��B�W��>�CA�qceO5{H�櫦����g�	|���#��
eW�0e?Zi6ƑM���	��Z�V��\����vmu�������lj7���lQGQ���u�L�s�%L�v-���&.*jI{_���,Y^�Z��YT��N�@��h��eH�����O���#^E��%��RCM�<H��R��9m1(�)�����F5TN��I�#ז����s���*"���-�.g�֒��V��|z�P!��:
�K!X���u��,#e��)
|��^�.0��J��xo�mk�3<�T��-Q�ѰL_�6\UX��225ڮ���h�õț8)8�j�ꄁ�ȳ7��d���JtŁ�qC	16�5��3��	z�ea�g���Q���X�HR��52];[��+�����q{��vT:�����rj�M�tzg!��5����nD�{.���(�[M��W��@��|�R��:�|��T����tӗ��iṇa��"����	�;v�����]��
k��Z���p��^K�.4<W��
<�8ӛw/4�4n���/�)��m�qUL��QR�v�5%��X֢�d���5Q/����v_�*L�D�z����/�����٨�p���U ��S�P�F�Nq� �k<��zd�,2$?i$3�5`�4=���I��G��`~��ʫ�*bJ\���[��%�D~:ɚǜ040�[��5R)_�0:��LC�ˣ7E�+������yn+p�4�8��/6��a�<���<~.��§�ᛂ��-�ݢ�:��e�	������1n��� ?ݰ�(��m���:��N,�f0��,�hy,���{�R@�>q�I���j�,b�Gcn�V������K�=�U�m�}����5�H���\���FZ��HU�
6[�}�k�Ā�~���a]k��k��
���N���7S�0i��)��ѐ��<�F`�(>��iѠ��I�)���b�X�P����d2��}����}�S��E������r��v=�������d�Zqf���҅I}Ս�Ar�K���W(g%s���W]�4�����[���������H��}��ވY5� �W��72K��F�<xD&�6z�7��.��ٌ$�HIo|,lR�=:�֝�O���'l����Ìe���b�ɲ>��z2*#��JԂ{�$��f|Ύ���+5q�;z��{��d�C3�œ��J���Q�2�댩���*p�������Fp��2����i
���Ƙ�t�
�(�&?���M�4���4 (` �0�>و���?Y&۞�-��B�̽"(�L��GaOqi�IpU�R�����B�
u���gD�|���$MK�S
,>��c[�p9��h�������L��l���"ŭMa�$�s��JB�ۍ���ƛ��!���b�u%���?}�TL�1aJ��N.�&��C��9k�<1o�G^��^������)0�>��J��TA�57S��UOJ���o������H��|&E���ۍ�8A�q kE%��4i~#�n	�%�Hm���IT9mej�JBaRj0�����{$p[���/F����ϑFV�h��z�XU-��v���c�]_�I��=n�6c���ħ��%^rqx�>��h�}���aW0���x+�jݮ#y3q���I���jd�����hi�>WeA���'�ν�`넬(�$�CrXF���c'�=��8�=�
��v�7��;m�3(�!ZQKz�9�(����Kw����Kč���Qߑ��S���B�o]�-��^�����qز����0_����R7� ~��7���/��2,d��]$����}x�#��㋒��o��O�F����ˀ$��&�@��d��3��O���y�^�ç����Sj����Q%;��O$'tNGJ �8L7�1�e�f��b.��T���00+Ym����������M#(��Lr�*֒l���4��z�U�_7�E�2��������|^<�B���*=S�����6R�7#�Bn�[��x�Q*_�5�t�h,xrחǋ�0g%�Q;���ͥ�Hr5m�P�%��=�0+�m��vt�5:F-�Q}4�q3I�>�^�̠S�Ǣ7jd3U_w�o@�te,����#�0�g:$�%����L\؉����61�y=�8Y�w��mt��)�B�ޣ��*%D��]�!T(�\���u�0�4��N.�pL�*҈c��v�ҁ����4�b���8��`3~��K���%̾0�d`/�2x���\d�<�ފ�j�>-B��c#�o(#��cwl.��#�����H⩆�z)��l�i��{#y� ;��P3K�g�o��ʏKӾK��#�u/�QK���~p�܀��E�jp�fr?L�^>t�}P���+_�Zr������kp����j�M��C�u^�b)����953r��cĪ4�	a|*Y�d���ID�P ��3�oS�n�@�� �z��JCw�!���y�Ӕf��f���l��Bch7b�x�O�e�Q;f�K��5��;�_��ӊ�I����+�;���"�R��tS`��q����BO���t��4�IQѣ&�h����qlG�"�I�{��~9��|Gf���L�����:����@Qs����$6<D}�Z�j�M�v�e��.�wMw���5L�	䎥m7I�*��� ��Hw�C�Ӊ3��hl+�m�*�˶r	�z��c���׹z��U�]�ܬK}R���;�Z��k��xc����8�64;wO�=+����)!���+��9[��^�"+�)8��TŚ�D�O�S�Q_uI��5:�B�$��#��L���=�<��
_!��tY-2��1��k�
3�)�(���*����F|� <4�K�ϙ�ʿ�����Y���IW�׺7�҂ϊ�"��`�o�^�μa���w�� �+�?�إh�h˒��J����.h�x�ׇ��QtlZKT��V�v<��LS(���qX5�I�}ڋ+z�$b�"+#�����&y~���x��4��J�����-�K��y��ťE�W	�]��ޒ��z��*��8J���6\(��6����t���m3����Zr�b�+ŋ������*�8p�	ܑ�޶"���e��γ��γ���;uW��)�?�H��[1���������z�;�jǨ��5�m�V~�Cj)�w���P��3�6�����{�����6�fp��"h�X��Ȑ�/u=�c~�B����u��?w�/�x�Vu��|��7N;��v�X+= �y��(��W,3�9i���ô�(D2Y��r�J�j���ɫs؁�t!t��ֆ%7/B̼;���^�V�`��,��F�mɄf�N�[���Yq<vW(ϯ����yv��8�.ݻj��Rۄ�?�-~c�}���-iޛZq�%��e�Y���߆��o-]"�^���@H���C^�7�ډ��E���$r� s�WA'�[5���1�q�D�tU�մ�Ԓ�/��}�,w��L�T\�5�Rc��-Rpv��&�"��K�P�7ס�2R�2�_�#�R��J<��L�P�Kb��F=�W���<�����q���SWA�ƽ���Zj_��
�&���jn�O'��(�"	(��`���Go��e	W����h��۴$��!�����T�!����)���3�� X�*��+Q�C�b�n���n6:jWQ2�ޠ��~�B*&H#'���Rśb����<U�����
��qݥ/*	-՛r�#R|F���²�	���ޛIb���,z�Vz���9+H�`@�g�b���8DG ����Z��Z�P iF����o��;�L<>Jl"{���u��/$�<�B����h�$�X���������D���Ҡ���r�22GV҄�N1dHu$.�Z�G��˾�5��L��B��d�h�*%n��.���(F�����^:���byt�4]� ��=��-y>x�>�� %p{�
�>�g���zcg[����2Y
$</���ׂ��Q��X�����q�u��>�3�b��Cϭ�{u����F1���q�b�
ȭ����m��-�A�R]j���Ֆ1��`wT=:���&���L,�zD������Ez�U��el�w���M���?aL�E��>N95=��͛�>����;�V�����,9�j�"��m�XL�9��ؿ��( |�Ѷ��}?J0mlŌ�"'|>�ON񂻂��2���6#��Xx��qw�(��2�N��b�������+";ȟ8��rw)_��4���**��YA��.S�=�?*h�"=�Cě�HX��wx��.��Z8�RM���i����A��:�,�z��-�t�>�
�$,0�[�������d�2G;�z=0��mt�L�2(�R�(����(� �F�c	�����\���,�es�`�A�ș�$�j�o�� ��V��Tk@�(8���yȠ[fUҚ��-�,��� �����]2�jp�᮳�I���|���p6Ü�	n��N�M4)����]1��}��)W�
Η�-���|���J�\`���Ԫ���^|�����W߄�)�_��d�ˌ8IQ}h�g�^��h�|:�AY��:�YTg�b._��"���ц�v��tx�"�c������W�
����}kl�ڰ�E�(E���'����W��܋���w��z���7r� ���I�w.��U$�$�M�jV�M�]�����6�j���@��&k�8����$hM�I��H�@�xט�'���Y�X��X;^nMOڲ����W.Q���,oL6��&�!��gĊ̼D�6���{a��ck�%��6NXL�Qyz������8Ir%�#����{���V�KmU�� HnP ̝�Ӻe���j�\���[���	��O�9����L�}$�w;|�K��l2+�,��ȅ@��;�{�?�
�	��7�wh0�s�M3��t��i�ʨT3����R����@�~���ʡz��J�C\���D� �Kb=V�1��7���0JT��2#��DS(�9f�w�^CA5)��Z���F����1��%�"uD�Yȥ5+�A4�k6����;<D��������FS�n���q*B��\	K}�G0���n�(9M�J��$\��I%h@���NV���	�A��K���H2y��Vu^���1b��W�[�'�]�xS���ld&��v�pᡆ���K��"���a6M���d��������|tM�`���R��\���q���c�!���r��NjH ���݊�����7��b.����;e��8(�/W�`����S��|;:�[g��V����2��D��A��`B�k�D �����}1~��hu�U��S��;c��H8G
r�w�&èNx�N�'ߤ�m�2�_� ��|m�5���]�Tǩ�NL���d��[�;2��0��!���Ы���Fb�o����'/^XG2�KQTB���Z(\�h?��g�&�J���4��D�/��-��ˆ.;5�ҏ���Y�%��ŷ�Z� �8�v<X��"67����`(�+�^�����.2�,���fqثr$4�b�F�a�C8����Zcm1��z�����J(]�9�*�h��_l�v��ƒȥl���7�zE�����:�\���Z4'�L��Fȧ z��v+��|���CU9����2�ܛ�ߟ�����5�y����.OU�*�
��יI��O�OI�5ͱ�,�Y�������Ec�D;ώ����e�P�Z;׆�L$r@�$��mL�<_P�����#��n�M��ؽ-|+I�7�tF�*�:<=��qN}c�b��ht���A������of̄�5D�<���r]��^���4՘�lv7�}��$�V��ʔ�{���1"�.����Y%{�h�ry�ťq�L�2���a�/� �"y/.c�S�bpe���,�Ѻ����>S�FVE��M6Gc=Kjx>B���M<����[|�%��ȴ{�[�DF�pDL����L?�R�i�� � �
jТN,�f� �I��(�5�9��$X^�� xvC��vF�5.ӯ�j�*ǳp6;�2�K����@��.#w�W��O~��Bg���F��@h$���1���l[�P��l���;�W��dוpYߞw�+����&B�V�A���c� h�s��:\����<�85�v��p�Y��<�Ax��S!9̻a�"�1��?�h�f[��J
��'!t���,Œ�@Cz����UQ�����~�J�H�k�Pi:񐃼I�_l����"i�x&�u��!m6��%�JgT#�������Ѝe��B�6���W�cX���?����?nzU(P���Y�0�����<t����+Ao�4^Rv3���
xH�4.���p�)_�5����}�L�>&��^��陷e����N�mL`��5��w|Q*��@Kw��I��Ȟ��X�]�È&^����g��ߑ�0����0�{Q�F8Jp;�,����Ü�X�8�6P�{�4��(\]ZJ��jo'� u��G.���a'���2�
C�=Lk�Tȝ[�"�\=;T�y���ު�x���,�blU���)m-v ,l�c��q��[��z�!'�Y�G[f�u?Dnw�cr�*�z6�ƽ� *�%�/�%����F}.�vcdW��l��3�5w�nylk�O\�����W]�#K5�� gk?�oL��`���
�Ik����-�ਏ~݋�`I0G���vj�[�_���+xQGk�
�q�	�)�vh��#ͷ��>���fp���N�֨�2*Y�T��u������d�߽�f�\��V�l��)ןk��v(���)��7t䎤��%��Q�,ƈ�9I0�F��㰳'k�܉�g��ī4��Q��,	a�|ږ�M�6��uB!�vҢ��1h��p�T-8#�P�ER�f�B%�	�4���6!��O�O� (��L�ZN��:zp���8�`�+B�P%J5��=���D �ԩS+���)����2���B�TG��K��|0��	O��bO3�⤍8z����l����[��e;fD|/h�[?/�F�a�Z��e��^)��;� B�vU[�1��cx@��<�L��:!K|s?'D��Rl�v����N�<Y0��Ͷ�x�u޿I³�YO�I)��j�Xe��dI�*�6���O%�ʹ#��uf~�_l0�ƅ�8��%4[}�\��_H1�;HN%��w��B��(�k���>P��|.ͥS�B��?'-U%�wܿ��B��]g�ɫ[$�� �Ura����S�נ��qo����0J��.�8V@,k�wB2����AYJ]��:�>������ş�%X��#́@FB9G
��ώ^\�r�x)Tw�jh\��%&�4���¶�C�9B-���Fbс!8 ��f��s��ۇ��+z@uw�bB� -�du*	/)�k�#i19�T��$�A�9N���K*�OZ%\N�{b�"w�j�y(56f��t�����R��-�o�H(�����1q7�	o�Mh�WJ�~�(I���ވ<��)�������
����Ị��Q����iE���>H�Ļ5Whl՜���"�l����*F�3��I�Z�o ��r2𙪤)>e����]J���KI��rh <\�E��Q�~���C�c8���Q��C+ ��ۮ��u�pl%��ETמ����Ȩ@ldt�sѪ���D�~Q~���'}d�)Y���>:�>�Rd���щ�jY����Dt�;>I�[?����ڰ'h��PD����W+�ٔ��[��. E2�J̀�QXK��h�Mo{N�ӵ҂���,C�!1��ю�AB�i�b�a�
���,����W�� CZ������I~�w�����+1lXc��AZ��u��֥�q4���=���^A{�q��~���3ܐ�v��E�>^��8�<�ө	������B��)zޒ?I��K��ڑTb�L����`|y�=Y���A�r�w�
r}�� e���[�_�CKV���dm�0����"�)�bvߣ<V�O+�D���h�Z<�$�����.���;|eK�F��ʕf�W�y?��`Q�LJ9_���v����*y�/� �-�I�1L�eުō����?����o�I�Htف�K�z5��c�E>х5��ϣK��$��������t��˛A��1=���W��Mr�B�cZr7v�BVߏ4?I��h3l9���U�&;��*�\����	oA޼�M�������ȵ0[�������<R�Q)�5�َ������xҰPx�I�<��_�6J�j�S���'5��_^[����D#
�N�Hx���i��������x���HaٷB�2��w(�ki�M�-d?Pv��~Ѳ�u%�iV�Y0���5�i����`�9,z/X7 �T�O�8\�h�ʪ��+��jH���CU�x�&�A@	qeE�٭3���S�~����q@)Z�� �}|�Fu��HӅ-��kWЦ����]���V��������sW I���xg�w�P2co0�+�[En>�%�u����Pn�G@2&"�լJ�㥻�� �A3$캷H��X�Ib���F+��j��7Ѐ�kih/�R
5|����H4��)��k���|�g�9��R͕8���ݞX�k���r�A��<��Z�T��S�)n�������tz.��p�{��a#:�;�[�	iK���>`�
̝K:��yچ�����L���Y��E���?ӣ�xb1�"ʳ��J{BE������<Yi؝̬VX"���7I�3s�n+�R�pd�#P�}"A��LZ$��ՑV10@�'�5���;,͐���?�>�F�Eg�Ea�t˪ ��'�T���1 Q����\q�SI�_� ��^	,���'�a1�;�Z�'r*ֈ�[����E��)�!���$�/=3h�f��P�K	��$s�%ר�H�b�����ɾ���+�����f��\�;C��eI��lo���&���a�����S�l{�j}S��w��h��P�&i8U�βc�!`pB�~-�B�����;��o����^F �X�1>� ����4?
�ۆ�:���x��xH�����oê�n���y9�4FY��)�=z"L�L��hF�kE����3�õF��
��Q�� �>mn5iW�7�G&��ϧY�թo�&ӴfC��l�k�|�r�`�(}Q�O*�e���v�����^�e^ݙ�.OU����
a��	Č���5�=c�h������O+���B��k7T@��22MeLo�KrS|�����֧���4X���:�aX��=�V�pJ��Wkmѭ�����`�P~WtN\G�t���NW�� (�l����������^M[V|�����w�߁���� L��������JK��VX�Zݧ�ӧ�{�'�ad��������=�~٘X_Q� �э�W�ڔ��=���ՓC���'Б��(�/��0�dA^��~���<�/�{a�!7���yj}���?,#�j�	���gpf��<K�_!�Q��3"<��z�3���2�c�4�ʚ�����Tُ���h� ��}�����1G��5��",e�[�
gP�a���=0�3żm�L���!���FS9[�+V�|O�Ȯ�-}B�5EDb�/�T��t�C�Uʐk�/bJ���Sm3�n���?�?\y����G��������ߍ�A��`lWN����]~sEG@;���Y2:�/�u�3--0�&Qg±�!�-�%�~eW�(��Tu�p�l��Ӄa���^C8֕\ՍYk��,Ǖ� ����2#[�6
����G0�`_N�Rf��$�F�oc(@u3C�/���.襏*d~մ�&��D�C�N���ݴ~9��B-��Kϗ��B*IT�;!¨���8�ܳ�E�G�˵�|���*w�����;���=�{�N"*��ըD�t���i���ZU!�t$<�Z��:��mG|0��)��t���;��
�0�I���@/�v\��b��M�mDw��1���O#��o�B�NF���4�ٟ�Q��f���/[H��Ϝ.�f�X�M��fLO�|�^�"�|�xIm,!Ԧ�C_��@ǝM3��u������5٢G�����r����@��'u+�ZA�)��y*_BjBsM��g�M9ڷJ�l��{���r�nϏ2`���(D_@��A(��C��C��doQ�ܩ��WЊR5f���<K����2y����YY���+�ң�����z���N�y�/���7lR}�� ذӒ����.xk3���O�s?��'��m�bz��u=��+&�f۾��6��K� �~��*u1Ͼm�R�
�`�m̏���m+ ����k��P��~���Ó�4��J=�g��uS��B1�����M������o�^u*(��"Y��m�Ra��S���6���F6x8�<��
�70��S	;	�0�)�W%�K���ۻ��3�?��y�6;7<��^)�J�V;͇�=2e���[eS*�����Q�sq����?�t�kYw�<OmWY.�I���Y_:T�$T��s>d���U��<�d����@�V���~](�%D�i�kCg�K������!}AF�6�g3߬ȅ�%�3�0ۭ�I_!��z�?�g�P9���z��{z��U���������N�ƍ��u����0��];��j(�)4�