��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��c����"3�t��%.S��T.K��8m0�Vy�[���
�����)rǮ�7w����اޗ�͖�_��D�-Q���
��	���DoI�4�{m�����NUc��0��ѓh��ǯ�5**xb��ŝ@����)Z���t�ߡ��y�!I��ulz�[�I�q�)�_�O��j�{�m@=��<WcZ��[��*C����^�����p�����.X��z�'�G����)�~n�1a`���靺��y��w��ȒW�T�1}�W#7b�~����8^��=J�����{�/i��5%Jg'!�rw���g�wu �P+}n���a�;�9N�I��ۚT�]M� �,$�шI�0Gz��)e5c�����R��E|�X���#R �ղQQ�����t�]˴æJL���1�o�x���D ^!���} s���ӣ$�E*F�~����a�k�{�v#���Ԭ� `�i¼�v�d��c�+��B'ir�7�ٞ�w! �zr���`"y5H�İ�G��&��f+&��'�Q�f��M���)ttm�$��NC�Q'�O�)�1Z�ˢEI�H�\!ߞ�g ҭtEuD��$$�ж��!���M{H�2��B�F��=־��#���V�~gI�3�},<�ѡ�=u�]�l��Gʩ�)��ͨ�`�%�y����\o����(E# �� ��g�B�U�?�����a�C���
y��I�sC�K �)��a�&Nx�P����*������5�C�`���B+��d�����u۠o[o��?�5R���^��@�+V�=i��7ڝ������,�Z��M����f��qF�t�<j�%U����T����#B���oj�Zil^��+F�
M.���>�y�ȝ����w$�s`�4{�JD�=���.�"rV38�
O�R���5�=�o���!C��Et�K�|΅����H�����
t��R���Go��e�DS����h�(�u��ufQ��n\��݄@��/UV�P��L��')����ɟ���m-G��M�
�-?P�)r�Z�m�x��N��j�Ő�������C��_�U=*��	H߸ʶ��e���Q���Nf�1;�u�{�Kq!V�ز���B��S���S�Ѓ�.'���6|�g5l|�WJ9��`! �"^Z�����6O3�-��x��u���~�q�4l#��%�d�O�.G������:NF}��򿕛�w�fꋘ��B���+��^��[����� e�ݢ4�==�/>K?����E��d4�w&���]�(�B5���ɞL3t��|:�a!���� �#*�>�s�ʎ����W�V����h�3\9�@nyR)v���L�.A��� �<�$	��% ~Pf�<�(X�r�>X���k�X�̡\h��ݖ�[G#6���H���;�����E/�4��!�O��D nK�n�wU��^��vJ)��/���$hW�,d��ȯ�p
�$�𛠬2E��h��׬[<���-')h�����[���w;*O����W�Iĸ�c�g�RKD�����vB�'��F� �I����=�Fu
f�3�A� ��H�(�!�fE���2z���~�|l7
L���*"�y
�r�Z�S+D��p��An^b � ��M�	 ��I$�Zč�7��Z���?<�}w���8��Rwi��?����pIꟆ	a;��y�ѤT1�j�(c ?4��LcG���G���:�0�P̓���P�#|��sd
�f��y�A��XJ�4�	l�#Z��b�|B�˫,T�
��_��� I�EQS`D����Д�y�:w{�S0�3Jet�ynL��
�KE�����{T�����`ނ��8������ϫ�~�g�kgJ��}���j�%�m�G}P��� 8�<���H-"����C���Ȑ�����vQ�n��R�[���x�\��zT��nd�&� �T�f</#����N�F=�ܩ��o�J���x�K9X�/
9 @�ƨV��ą���N�e�T4��vM������Ȃ�A�vג�o�+oh�̉��Clv�m�_��13_�C���.��1P�g�#�q�RH�+"*n���*~�^ ϵw����-����,���/�0���k�m�W�UZe���C�}��+h<^vѸ\�:_�}�A��G��&vO�2��������(E��
v�z7�������0x�F��G��B����tG@I�mM�nW�0<����DA�P�Fw� &/B:�
��(�9* �X]|H8�&���`SՍ�톈`�H�k1�9��R��no�L���d�C9�n�A�pL0�����Jf#8	�S�_���'I�O�:t�S;��ʋ�m�N _�=��m��.T�T )M���,�)Y[�t��;Ь�!Zs��`}�q�YT�Oz�\Bd�%HՃʡ7�,������~���ೞ��o�sN��9P���6���������X�j��$�� �<)�K��j%Qt�VF3M��_~Y�,�{]0�0��k��IA��x����fڕ�����x��"��8~+-q��='��N8&&C�
a�2�;�N s ���!�+ɏ��~�~��������KP��v�u�6�T6���s��0i0r���y�;"68��_��_���G�L�Ra9%�6g���Y��{�z��C�0�c{�P����l%be�#�^�@r�Jn|���{��kD�$��cج���e����/��p���q���ױ�"�S�D��%S�]���')�+UT7�z���y�'1���"ӑYτ�d�(9aCƜ�6Iq�/�	-ғv@7P������נ]{���D�˜.dg����>�V�&'���������
������b^R��٤����'ߑ_��=O�!���4�Ԙ�w��n�c-�!G��I����w�ś�L��6���}n�u�{}ye\��Y�?�ڝ��"��ތ9>}���Ŕ�G oوpca��-p���B�6Z���O#�OGf ;��2�It��o�=�ܙL�U`���Z�6��	D� �򐁁���#*zCK~� ���� MR�D�ΒUm�,^�p�2��2)e��)�2��K��:����\���p�����}ͱ���ҁ��ĦA��a�t%���Ej\��U%��ˍ�z��޳�����g�ť����;&qf%���s�B���o�}CB9�NI��2��j�r�_�`�ޜ�)&
٨`b�up!��?������KjT�iX8�`L�Rh_�GH�]�Ӳ�� ��q�ò9���N���4��*Rf�7	k��ߢp���G:�Z+��8�[X,a��tĳ����}�}F�y�Q((-�����;�Q$��W�.rh�ֻ�:n���Q�4
}7m*Ix�ak�S���X�Z�,��G8:�_�ƆrO��Ĩ�Nr����]X��E��[��E5��@B1����1d��ND�h��5ov#Z�x|���確�C�*�sA�u��Ĕ��vV;g��e;�ܾMK������p� ���r��SƢ�گ�&�4rT�Q���Z�������kyr=ٳ�֟T���<{t�],�W�CןL��/;-�\���fYZ�>n�j�{�uXc�)�`�b;}�<��d�8��k�����5�MkK�P�>&�ӷ�߭�[ZV�����}$�	ݏe�9� �j#�j5hE��qE���p��p��R��_���4)�АPʈ5�Y�0�p;���<�{�7�j6E�4ڰN�Ye�=������W��j!�=�N)��G�$����W�=[?�j�>��I6��+k��Q�����ۨ\jܩ�_�-��nd���)�Y��;��%�ǲ.J����.����V��P����������a�	<2S�#'���a+����ýM4�m"�t�\����!� I�TzeΝ�
׸��.V����В�l�	����T�����D+c5���� ����{����\P[?����ND��Ԓ��
;��Ѕ~�h��N�)�: �$#�N ����O�<Vu2�h1���+�4{�nИ	��ǃz�8��#;:
as|�2ӕ43�͐�΂{�P��)�-���B�ƿ�Jk<��_t��6�=;�ó�ѳ�s3�;7�.�)�ؓ<�Pm���d��RB���N��L紡	+F�O�	���n���X߯9����P�.�t{ʅ(\u;�Z��ǒNWȠ��}2p�#�)�U�V�C��25���wOٺ���`����$�D����*��� �W���q{ft�T����zp�o\9����Xe]�(��zf�[��'�����Ml�c��whP��N}&.1,йYy>��r�����a�j������NhA�Sⶊ�*0`���� ��W`�'f3�O0�Kz.$Lտ`� $P�r��g���L���µ������dv��쓆�����(`U3���ʖe ��wR��  ���=�H�~���M�x����
�2��,�8G�6cP06��v0�#��+vRl�υ��4h!(%�@�Qi��-���ۄ�ٽ	^ uΏm���c+-$e�j$����ݾ��~��^���s��vb�R(.�.��2o.��z��F{��w��ɋ�9���7�Ў�6)I1���?�ژH1/[����������湉~ѽ������F���ǰ3d��Y2�:|��&���s%���, ܼ���{�� ~��i�f�c:�U���$��q�h2���\G��%�o��<���&���^��D�5=P���=;��oNݹ���}A_��N��I��dm������Ám�fW�v)�������p;i�#��������F�t4I��f&t��p����ux�=Q�xs�X�i��ڭco�����u����Cܚ�֨
��{��x�>�w㨞��z�j�?�X$;�q�A�{��;k�¸����fSWwn;`+���6�ڀa�q��.�K��c��@}՗���a}~
^������k?>���������u>يI���ػ�B��݉�'[+7�؉��
V�*�*EM���6��iZ��pFՇ~�r����	�����@����W�D���O�}��<�_o�%��(�d�� ��+�<dy��PX��z��=�O���S�y�1��h�
GJjlb�e���	]��9$��,��ɉVf�y}�)����ؘPЦ�U*��JEw1���RG��ŬD�`2PnS:�<}�i�M6{�_s9h{���[R�9&}��8]2Ɋ���Tȑ_J,$H��CE&�IZ�rHG�;�.��#l��t�/��dȿA�AgB�D���"g��?���"Z�jgn�N 
&H'���iAm�զ�&<��b6����v�h$����'&,�d�L^�E�_�C���sJ�/��Z 5���
8�j��8P�Vm�"�
��Y�[�%Z�g�t@�ă���ď���{�84ޝ�1�jK�{b.,�Y%�K�!}/�y]������Pn}�������I���bi'_��q���$;�lo�t�%�DK�DIY���/���ͪ�]9���lf��x�W-J�)��W�UaTrb�U���-W��y5�ٺ����hFF��9�1��d�ϊKe��X?}٣�;��x����"���@*?�t%s���-j�@�P��}�tL&DES@��+��4"�&�a�1��ɻT�����(hP%�g��a4�t4&�uG��(�c^@z݋q%Ȳ[s�@��]t�+^�\�jn���JG�c�$������j�M���V�f�Tz3����{t��{_��_}vf3���&�:�%'-JB��~u�0�&�л/׉'Ϋ���5h��b#p����������f���[� ���nkIc��x�X�ǽ���i���9��lD��\�6��y�x���{�D-�J�O�Y*D��I,=���Ӗ�.9Z��_iue��Fb(B��}��`2+P�N�y�B)�4��C�W&p�6���������ulG�� ��j���~�y�TJ���d�Xw"0�
��JG�0l�fD����3<Bw��iC�r!M܋b�����ZF���K� �<�t��X���?�u����{t!��!�
�fo
/;4�Q:,O�k�T�.3%�ۊɟ�W�ՙ0��N�z��\3��%F1��i�#��]�����.X�l9����Jn!jP�<����h���;�c�����(I�Y�gl��A=D+�:Љ� �*E_㭚�SO���!)����řKp㌸�U��D�{��7�U��Ȭ�a�C_ᥳ>�������U�@	t���|S@ź��>��1˼�ow���IA=U����́2p�9k+]��#��Q�Z%O噥_|�r���훠%�ǜ��~�[~cy�vn��9�4�2}��W�B�|��=�s��C01kÕ������(/E|�\4߾;���V�cԦ{DѝG�|�z��c�R�h���&�'��!������^�I&���/$��Yag�a%2��T��!����_�<xEI;!�˟�`X�p�8ݑjY��{*8�"�^U}7�Y��R-�
ҩ�'�����H`mcOd�O�̊yB�l� ��ǿ�.�=Q�J�2{]%�5>B���c��g�p�� ��C��L�LgӨvOO�@���P����Z	��o���Y^�1�*n�ʂ�l�vp�on1�YXq�|VV���~>�x�%eƵ��a��
;���ʟڹ���A�V�|��Q{B�0a�]�j�k���'VAtf����C�7�.�q�^�k�m�u���@��H�pn�D��X=A_���B(�8�_Q���̤Q���2�=�U�?!H�`!�X�7�zx�X�7V��=��x#G��1�����D^
�m۹����h$߆��e����t�Toiq.�����rb��M�Uº�����|�.��'$���%[�N:ݡ���U߄�L�8UF�\|,W=	O���ϝ����!v*׎
G~����<����VB����K��:
M���������D�{v U4��7�!i����WOc�Xέ�?E7�Ap��<z
�����'O�4Xt/]�����쐉e������24/��z���22W���y=��kB�A��~!��
eZp�߽/پ�HY�f�c��bNЩ͠A5�!�rv2���=�J�aN���ݣu���s䨧�ZO����3^�sb�E�"��?Yw<�nOG�|$���^����z��y]�	��ŏ/��R���E
U��&P�C<}��zZ���� ���e5����K2<%ؗ�`i��� ��7ǳ��`���w����GI���_kx��_�(�J�|�m��m&N�vi�8�}��U2E���B/�%9ئ�:F҃
=yZ2oLHV�f7�$^DB�'/����yɕ�or����қp�ƉA����X�u�w����� �
@�v��W�?8KYB����9�2�ܨ5}���8T�6�z&�$�e���Y���{�5@SC�f0��Zd%bR��sۜt7.1�%��I�I���E}*�s��SyH�>I���T��r��Qi4���u
.���x��0emHU������q�I	�L5S��C�Q�'Ix�x��G���dmձ�r�J�n�$T�c�Wb/ٻ�'cPcD���˚�J�r/f'lXM5�p��=X�e��j�����1�FY7��t�s��h�jM�q���u,��j�J�{����<K?����uc^e�w�*�-:f\��#Z���S�&"~z�<���۬���
���9��>>S�2�%��biu��P{�U�	Z����F�䥵^Ϭu���@[x6�`��(�4t!� I�5�Mp���i/	���ʸ�9�3n4*�����6�n��mm(|!�4V"0��t�'DE�������{�  �qǷӟ���FOy���ۜ ����t����)T��S	��:�Z��j_�Ȇ������s��k��҇�Ȑ�=�a�c۞�����I�n�ݤ};�J.�d�w�mW:��ut�����ácC(c�j�i'�)�KS(s22*�'�A�^�sz8�oS���;�a�;99IkC���=��,�@���D���E}��#o{Ʀ��M��4v>�4�P,wM�Q��:>*��5�DF[��v�$o��+K`�N�]�Xx%~1�Ri!�k�OS/�665��K r.a*W��{��ڵ�N�{\{ӹV��})���ʐ���Fa��j�æ�n�Ad�g	ML����#˾uh�L X�lYJ�?X�6Ry�0A�
E}�OX-�����.x��9������M���Ř�If~�����7j�z�`rĢ /��=��>�'"��R��b]��x�~6�����v��.<v3ƥ��Š�j_�˾{ڙ-0��85f?݃���B�Qm��X�9�z�U|	��B���T�A's�?q<.Ԣ{��v4KE����{!�в,f��H	o�kKs�Qr�3Β�=��v��S�M��] ��@~˒b5;��=k�m�jP)�?�/��NJ��&��Ul�g��8�ҹ�[Y�u3QB��B,sEZ'��G'�c�?��2i<V��%��:�����SшG���^U��#$�G-�
=ea)\�5��e�[�_wktc�شvИ��?\W|	q!�Pe�?�͊>�O��$>�:M�c%��:���i����[��r��*>��}83�w��L*��v�,�E��^�*N<��̀��0�c���Ĵ���8t��+�\l]�X\�d+2�#��7�>�f[�юl�i��*f-�*�!���q�5�b��$�)�V��0}<�_Y�5����0�����C���+N���iU>\J�f�vc��1^�T$��S����4�����:AP������v�v���g^�Rk)^T���gN�2<�����@G�����,4G�^���C$����g#)ѹ�v�#�Z/�1e@��w��a��e�I�*��K�KDn�e�]�F�Ƈ4�jGfv�зsu*�/�Xf�0����~b�#�=]����L~� j�A���e{���<͌��ǥQ�lS�Ѣ�}-��-R��7yTy�\���.���=)�ǹ�J�z��wI�-D�񄝨�,�2�-��dnA��SY=�8�aef�,M��A}y��5!,��x����aT*-��A�׊��i��l�՜����q
7�q~0L�܋�8�w��v�l8X�wZÖ{�thc[�Oi�ɫ4���5w�����0��SE4OYDE�/��9s�oE����L4�Z!`���E\0V�!n�����ܛs�k��'6S�M��eJ�L��`�4s@d���8�*T��k��X��\������a���	w���i�<���S���t]~UNS�pc��wƘ�+�?�r�A�hE�W�W���S%�
��>�_A���Jf�3>N���&���� 7=Q�*Ϛ,��_~�?����-D�;t���,���8��]�Z8�~��x�w!�*����2F����Bb��͍0J���C���bQ�,2�� *
�e��Ѥ��:�G9�\O�%�i%{
�*o��1m+v�M��ˈ�6@����6j��iK�Z-�vM�p�ʽ��7>�&h� �Tk&�#r�u{S�붿�7��L�M�]�#���e3��xU�hf���_~���D�6S��ٍ�2��|;3��Vqk�nL�u���N;߈�Ā���&���qa+��k0в��7S�S:��<�t5F��0��^SkN"F�>��q�~�J��!`z�6������!)�=�Vn
�g��� ���	`�;���+��S������ĝ�ɩm,�A��a�$��e�&�׉�=%�X�;��V���J��֤s�h�sQ	s�����_���mA`IdW�$�\Qι�%�m��j�v���ʫi�2j$=++���&�t�����d-�ds$�
���݄&/�:5��r�oUc�W��ɱ�+����)W���l�^+aM�@�D��+���;B����j�l���3�X�>��Xe�y���e���p��u:��;ۼ!��]��(�dn�*�<B����Z|8HH�s��Uf6/��<I-�L�e"�V8�8@��3ĉ^�HH�or��O!�#;�h�4D%���G���3qAP�&�w�"a���ܡӝn0��������>�L�U��8�ǈ������zE��,�7�f�M�Y%��G���_d1�X,���c��F��7+(�a6�/��+����ʎo����{���,�����2i������G���ن��)�
W��|��T���o�\$~���{��?YR���.yMW��@�%���������ʟA'�شk^ ~r��I�-*Xs�T`��=�d4���EFVȼ�3���ӇO�h�����*���º�E'�sKC�t��,?UΤ�W�Q;]�,���O#ϨzG��{v����$��TH�o��$k7\y}*�*.�p����χ��\��������Q7v��a ��JXqU9:�[@"���>3pI=}�]����y�5.��&��Dn�h��9?pe�Oٗ�h)e�c�F	��v,�t�Z��񭛬P�<pAK^F�1A�1���JV��*��"��k�$-�ﶠ�%��a�%O��\]�ʛ[Kw)(\�B{����7x�U|�!^����?g������1N�9`�;q�Vr��T�Fn%���kK��Q����@��I�;��\��p�-J�U��ԇ���j�f�i���C��$�'���X������qȽ���]��҂c��}�{?�"��2sG�[���)W��yz�d-�j$ԣ�����������!uemP�%�J[k�K�����cW:� �K��u2�jj�38��\��ϫ��ш�rM��k/��)��ROA�o�Q=�Q	�KMmTk��c�}�R��ǥ�:���ύ�Ѫ����0�k�ɰ]���o��L���E�K��h-29�C_���y��AZ�v�/%�%��d�뮃T����#H�9*=�ޞ���8Zd��9�Q���ck(�v5t1�.`�uuH$3�l�f7�u���HֺjΑ��n tm"��nx �/�:�jTR�:a`�;~�̪��\��x@
(��Z�����:��^}<���R��.���p�6�zu��P����=(��?Q�R���!%�ך�b��_.u���g��+0(��c���hp�%T9�.�[��C�2mX�����^����]e�|pƼ��Z� )u$���^t��Xm��+nֳ�N&��Vd[�?��L�:f�Vqt��sсh��4;\��"�����+ZwN�����U�}��8:���Ub@���g�cN��ўĸ�vU9Eyú��8+ H$8:��Ӕ��*�l�ݢ��,�<�)��ɲ"~O�ƙ�#���:{L2K�� ��yZtu�=fW� ��A�H����	P7��s
;��;���p7:�F�m嶢�Y��]J]�	�1�U�p5A$H�"F��Z|�;b���L�_N�|\[��lEg�����C�۴���y���s�k��Q�u?0�٫(��q\m�G׳}��!�;��)
ܻl�tW�$1��T��d�
3 P6#�9�=���\
�zqk,%��S�$]�H� �5m֝��ߣ�$V�x#����6���b4:>Y��m�Am�����_�zfx��$�� �B��I��G��I��&rrt:��]㢖��)��5On��Ay���O�+U{O2!W '��t�^�j^�����ט*)�f��Ҍ]ws���7U%�Fl���C�;�*	�t�Sn?{��T���JN�YM8V�_Y#��s8�k[�?�D�
f�Y@c��o >��p�\�ߧ��/��WL��udŇ�-QĒ��BD�D�Z�,
Q!����8�d�#9�Θ#�����6z����Ճ��	�{��^�\3c!MnW kӁ�h�p��}�+Y��`����2��l��V���3=�#>ͼ�T�*G�yޕV�Y@��k'1�<W��6#@IJ���;7a���=��z3��.�ue�y-�b���,��硫��X�'�0�}�srҘ�����ƂC�#ј���}�c/��}��>��}��
~�+�l,|��t:�BD��푓� �j�_�6����\�/�Ν]�g� @�D��7��.d�7-_�sG62�Q�t�ǌ{��nU�7�W[�9 W�Ä��,TL3.�K���+�;�!j&	��|��+�K�M�1���'�9��թ,�M��2W�/�k�p��#|#�?I��*>��$ɟ���blɟ5�N<z�b�I�xKA>=u��W����E6_�A�E@���Ѓ��9�>C�_��FT�������u��F��.�"���Ȅ���򦒇R�e���;2�O�+M]f��?eO�צ�q�s)5*�nj�$��`���_B�(�i��&�ڼ������%�B�L�RRT�F�޿y0�<�_dA�}[e�i!|9
�r���L*~^�꾽Q��7ܽ����zܻ0�5x,��+�|�K��=���D������?���0R���a�G[շөY���W�y���o�7�������a�IVAQ���$P�`��iE��n�z�R��R�DpS{�:�7ȇT��M'�[B�e�0tf�F击8Δ�����O�H�P��ޢ�$�¬�tTHM!��1�2"������&|��f�-�K�{V���N�՞뢤�-�q�B��%�j��!��q6�g���o	M9/��݌M��wY=��j�g
���9�{3峤E�|�~�)�_^�LSr��Q3.�V��3����_�(���9�-���q�K�lm������J\1-���xz�QjR���VJؽ����d �l��Uu1TG.���p0ѹx��b-(�.����C��.�6��
���.�"z���.�7����0}�g�g�5�X��(����䟉X����9xgF6�@�c���޶@眚�����HQo\^�胛?�'c��םt1ꖝ�l�,*�s�]*� F�!Ϳ���(sT�ջD��E�_�$�B,w�G=ר�4���M�@v�.���"n��
)��B-��)<e�/��|Y��6�$>`�3�ƥUw�>T����5h~�5���>VI�-�z2 5��u��cL�xq�<�[ ԵOB��ٺ��ݖ�����N�ˊ�jN_��U5��ǽ��<����mw�����dX���:��`0�?�S#B
6ܾ�i�B^#�͜դwK�!U˦��9�?��<^��-�r�v9�t���
�B=:D��:Y�c�v�˳N!��\sD3����B���4p[��b��t;�v��<1?،����m����Z�A�JO���Rc��FU��z4]_��Ӟo'�ލT���V�,I�w�Wk|U�<���V�5�]��/��F��~q�S����k��r�0�<�^��	��O�������/��-֪-1�uf�^�PwC�x�����q����wz���G��Xz	D�{��R�׉��KN�}���E
�q���t;,��#J�2d٧p��2�Pi�Z� OL�m����z���|�����)�aB���D���e� �(�}c ��J��c%�F�2�Í�� ��:Q�On]x�v��W��r��^*pWe=ݣ7b%d�#��F��#�|~�e�F��_�t����"T",��v��e�{ ��jiE�O(���;�W��Rj%�U5��M������L��fܢ�ɲ��/+�X�y��(�����$�6�5��FqP�Y>�mU�ϼ����a6RsI�(U>�
r~�P �S�T�I#:tT���/���)Y����q#p�z>���R<c��!�ݮ#|eML �k�h��i�ҵ�٭�A�5�Y��
;a]�8ͦ4�_��Z�ܘͣ�Hi+�vE�o��h�`r�c��މ���t^h>�G�est!�fS�F�����<8)]O¨���6��5���>8F~�aR�\��k�5�h�Y>�̕��y2�d6t���m�a ��>���=��?Q�/����$�<���#�+����?����6����4����DD��Z4~���#�;��O��A/ǚJ쓺��a?h���QD(�
�M"G��~P�0� fH���J�d4�!%i�шK[���/doh!��2��SC	����#J�^�չ����B��JH-%�}��58m�rK�1^1�u'\���Z�q�>3!3}O�>|���UeJ��B�����;ކ)CP��|t&��;����:+K�W��~�Z�i& zm�^nS��>t�/�&?���LD֐�x7v������m?6�m��.E��L^+�n��a�շFr�N#|�/d�!�
p�D�>B?�����e�F������b��Ų�GX���8ًYr�!�X�g�F��9Ү?�['��W��O`��HmV�g����CL���Ì;��+����f��!	���U�'�� �Zw���30}��i��+UP�b�*�ἅ(.���>O�Z�������;Ŷz��e]AҎ���,�g��u�L���4.�Z[3�n�4�f�斚c\��	r������E/y��2�hrO]���;���܁k֢I���^p O/��f��a6|C4���n��
R���ߐ�0ͣc��Kt��p.esur'U��(q�M\�0a��a�7���[�Q���P��K��pH"Գ�]P/�Q�b	���r��2 ���۫v1T�Yq����)���**2ފ���s��]�V��.��r{';��D��v�9�[&��֬��lM�:��i�bax�3�II}G�8�H�K�#������x���
M�@x�D�a�����V�z��V�,��}e�����@���(?�\�⋃�W�S�軌&:@�Ɗ�Ls�Etj@P�mb�(S.������^!��z��3���ah�~�(p�9���a&!�F��t6�T��O^|es���ZشKG�`M�j��l���,6NLFQkX�(W�l}�	=U�1�Ńڒa=�>��IS[4K��S.=8�ȹ,��^@�zY�� �VT,۔[W�<�h�Rol��7iQf�0b�Փ�~��ҤFAs�w�]��s���k�*�^�4ù���qNj{��FZ�K�,Cѷ����G��	&��Մq�4A��w�q�
<\��գ2p(�9S��O81��0�
��u���od�ݯ >s@Vc�#���^m�$9�$"ǧmw�ѧ�5�Q��W�U�Y^�k:/G~_*6[����9���)�:���ʩ�2*�sĶ%��M�F����Q8�!����!tv����ԩ�2K^ ���yZ��	�m�z4���Ht�������%�)"E�/#f�kF��>��	�g�5�D�f0�0p.�
Gր~h#�@�@�߁�d�җ>�#|RA�v^�W8�X#�2�0J,X�|�͓��.�7�<4_�Qm"����A��{�LPU�K5�]W�s%��!��R�m並��R%�K1�{��� �]^�~�ç�9�����M{W3��5u�)XZ�ո�nFDHt�qD��6	����0�������N���/���]�,�&����r��:��	�q�֔{&���EZ0�^Vl5�����(�_�����`�"�c<�� ��i֟2B?	��[�T��7
�zj��)��P,(Y�e�vI�u�nu�*�y����FJb�fn�.� ��9�<Y	:N1��8[�~$s���7���s3[�@s���W���jk�U�_p�#�������D�*s�t�aZ�&�7��W;��@HND!s:R'�z	H4�#�"-9U@$J>�E<B��{�{�6N���/�ǔ��7�f�	7� ��(��M,�`��Ԇ��B6��5��}eȘ�W�55��;�$GUR��M��"�'%���+L:����	0��2��������k��[ŻT��Z��#���z�����Ш2��	�	uo�`�UZt
mRIoΪG�:K��a|ק�pTL
)�>�k��Y�5��NEۙ���%Q7 ����^�N(�H���.`Ǜ�jӯ9O�G!-�Ë��_^�;C}�sZ��-L���q���v�����݁�	��dҠ�����0���%���LPqe=�D�|!�7_6����`�}z:w��7:IѵA�O�Vw���1���V}K�Ư���
`�f�7��K!f Q,�$�|r`Z�N�P?^$��W���f�T�PP=wf�! ��-��a���(�NW����T� �=�Q����|ۆ�/�|�h�cQ�HQ8~夽 SW33ܱK�n�8����0i�NH��,^%*8���0%ٝC���.����ƫ���&ݽV����3��X�Q�%KtG舗݈�@�*��!f/�� 4 9���L��`3Y7�	�7��8n�N��jw�`L�e�Oe�Qm�ԝ��r�W��]6@���Xt�yT����L��(�#�K:z�"�W
=��1���Q)"v#[)~���q�\�J����H��GE����$��Jbb�T���@�l�z���+b^��:��S�+��a@;[/�|�[��@��I��^�`��?��x����Ӷ�}~_���͢qo<]{���u^�����W�˷h@O��rj�aQ!ݿ���.XMG�i������0T��E��/<T�&w��S�-���"�lS��o!����2�B���kl�H+�N�d���&�$�̴�d�G0�&����-�i����x�G�˺��0�Go�+��y��B%��d�[�L��iPV�Y͓��_\��R�NT��:x`�j�#�ƴ,������*H�^\��o��9Y���m��L��W��j H�����}��p�HXX;�ً�L0Թ�zM�r�� �;��װ��)��%B��ו0(f�l���Yn����ˡ�|��X����ʫռ3\}�����'):4gY�JC+������I�z��7��e�^��$=�wV�dc�1��W�.\^.K/pGk��,�t)��z���#U&�W��KV��EZ�%ؐjX�*�����"��K��p%�_��C�S/�P���=��9nwԤ��V���a�q��bl��u ���T��[��a��qJ��{�J�-�",9{��G�}�M�<���n�*�q�}^�M
G<����r���_4�2�h�a01��������y�%N�Z`�a������%w�b�_v\��8Ks�(y�]�h�B*T5�j�b4�,��w7g�j����2�X(�Ϸ���)�$���\v^���W��@����W�[�d����B��C7�ҭ���� oċ�:HHi*M�p�,����D�8� ;��Z����F�D���A[>U���M�ĖR��~h`j�0��R�BE�-%��]��W���r�O,2/�Ǚ_8 �^21�v���c���%��G���\�dO#���p��d�p9 �@э���x�#��s�O��Eg�쉺'��8x�d�Y��To���Dg�9Jn�h��U�c��@�$}>R.��٤�4H�RK��H������f���0����1o�����������=�&?��~΃Ϊ����~g�d��|���K����Y� IFŐ��ڴ #�M��xֈv�Y
���@��@C;��~�QA�0l�gRE���O�Яa��o$�0�{��%��ސh�2g;���,sͦ2
V�/��<�=J<�O=��� X�f��!L$���7�/7�}�>��f_r-_�'�0���X�#�)1p4ڹm�n���-��&t��z�,��Ҋйu�գ|��alh]�a-���a[x�M��8h�5'�!潑W �ŝ>5 #��X���j�]�e,<r�Y,SE�z��\��_��"��B�vd���P� �-�H���tN�5�4�˭IL<��Po7���M�����L秹1�{�2ۓ�̑�u��rm�|3���˶�x�.�]2j��x���H~�p�׊c��Zp�pp��L�H��ϫ�x$x��D�L����vD��:;s�
>�>qs�R��ǼfI ���S/b��.��Be}�4�C�C�.� �,���W�<!.�6�)�[�I�F�i��3���5_�i\�UY����q���N(2���~�"ZȻB����ib*�"~V5�qT�߷qs�5{�R�ն���z�r�@�C�P��� �Κ�Q�a'/�b�H���[���]?
t���`:D�
��br�vKf�;f�lvSjY�nG4�?91�'3��rK
�4ʻ�P�I��兀�5�%�n��,'Dܫ��i��"!Y����ݐ�X�<�1���&���o��+��xJ��:�V��U.�~R���U��O��5��Mu�x�K.sz��D<���B
���L����)�e�W�)N��!�1�棷���t�;X�T/5�a4_��Ey�/�$����6�-��C�[�m�.}��4t�xOt���s`tJ�R��M��ՁTEn�&7��-l���](��kc�2��ę[͙W����C�B�Ph>��3�	ܵ�������fA��iÌ��q(�G��J�i��Q/��/���8�분�
}qp��#����|���m2\�EBA���}��_�$���'����jW���Ja�����%+��n4㢣�<^VW7�:���Z�+���;c��Y~���:!0{�uG�����E*3��ӷ,�f�9u�=8�z}� �-J����n��p�N��WG�͊�8.�QOf~G$����[�y����S8JA���I�Fjd�pJp!v�t;�.��_JNk���	̦k�g��U~��ޕ�O�e��u�h�E��$�پ�M�
fz��"��n��
:��z�Xғ�{���}	uH�*�XiO%�Ď�n�a%�3=�,���N���Q��?�pk����)��;5�P��ߋ�2�LC�Sҟ"�@�D��Z�/�?��̓��yQAX�ź&^�~�#�x�*�䋙&&���Q�j���~ޔ#���wrG���H��TY��
%�n�Z��� ����D�6�Lm�	}�z#2~=��O�m�8𙝽;wf�3yR+ ��ϰ*�Lt�O�[��,�r�1�a�����ߺ���D�?�u],�a�+0���̷�M?l��UA�I�<g�g ����SR��z5�z}?ξ<n�]F\�C\Y��	ƣ𖱄�M����/���y󑑬���8�2.u�L����%��qt�$������0���j�r5�����������>�<�]#]ˀ(ް�TI��0N�&��H�d�$w���n9a燿ի���t����
	_r^#��4�ڈ� Y��0x��j����ѥ^��z�w����`�(5c׸Ȼ��1�-���{Ug*2�# �z�bz��k�g��o���.<�Ցi{����u/3�1��p6ǻ��6��F����4�	^���[�U����8�L[��{^��K����e�"z���b	X9-�jc��e��]cK>�%Pn3��x[��(�U��Z�bš�VE��;�����>��-p�������X����Z )�[US���qj���ч C �6�hp~'��޳lW����������S `�Iqٶ��%>4:�L���2�-+2M#�vȳ.lA�-���_��2G���b���Ya�L�p�:��z"��V�+��vd��[ b�9�*�-�sXU:�k���4-�o��C�J�k��J��q\L:L.����H��Zga���=jfI��)���ߐ��Lsu�£ޢ�5�iWTBM���V�5_T{��IluH�U��z]�����D�^.���E��/i�J3�Z�J����aN��Ʀ��d�,�	nr�y$�D�����^���>��y�jc��b�ڃ�"�'�=�$�����#�T
����8��g�����bəI�2��e����@���4%��;u�n�A/2֗ϡ�}1m5�lJ�dT�z��1T�"�a�{����s�|Qm�h���[��t~�f�X&��h��`�-���<���5�jxrwIծO&�e�-���u��&��/-��$�+�2R�x����S��l^+�����U�
al�ъ�r�7(��ap��v�U�vө�:�B�f�k��3:Y�%�4�-�?U�y�����Ǐ�q��`@�Ay˲g�$I�����~����0X�S�eR�u�����5[�,I�ׯׇu��߾��zsӒ/��Op�����y�����}hM&���ؾ"t;�����L3�tL"9n.r!�|3>�B�g2��>�d4,`�>���c
��#��t�&�m~���/g����A���G(HeM���dC�Ng',�[\X��qKG"!8��]Mr��� LL І���ːF��ɭ��Ĉ{�k��n@�zbD��ךΦ�
1YW}B���{5�\��o��Ȱ��
)��o�`^����A��=*��:`ף75�r���hՌ2e��R&���,�]#8ȡ���K�k���/)�S��NW�[����"�����r��>x9��(%3�/�,/��U�In�@�p���l�<uW��w����@��o�������χ6���h�g�me��}�xכ8��:
��������U��j�8�ʲ��j�9(�{i��r
A�'���޳\}2�15���J���st|�Y������#�@~G�&�3�����
���w��0���L��խȞ��O,۶Ш}/��܅^�^�>�V����	}��!g��ډڨ�YQk�L���6ŭ��H�0�?>4�1
,zǙP�Rd�����߹�W9�Ss<��J qR�蔞4�x�5�0Ea��Vh,:T�nl�Ox�DT�{b5{q��秶��nL+�b>KH�Ȍ{����0�	�?�jb�����r6û$���MGFX|����py~��"�fH'�~k���E<���3����~���ԡi�[�����ջ�ܢ}HT{O����CѠS����N�N;nl�0<v8$������vk�s$�ꨄZ��%< �z���u��}��o�齬�-@��9z�@�Y1�����\�Ahc�P�S[P�*�(��x��{�t#��/��ܜȍ��Q?�
b��@�8����=3��4�74����2�'̕S�*,��Dt-�T�� ��x�ô=�p���?p���ia?\�O��^u��z�a�|���懲�HW�`��e̩��GjWQ* �^R��
ґ��ۉh�0���)��X�`+�)���]W6}�
���h.5��'N�.�jZ��uYe�t�.��M�g��t濧 ~]��5���AO�;������ݡ��������/�?'����<r�x��w֫gӱ�;9�K@���_9�mx=:��3�+տ'��n�̜�_޹㢸�>8�u��bȧ��,���wSD�ڧ±$�c�c�75�^JU:,+q	�(<�y�XᙿTN�x��ԭ�u̕�k�W�ɬ��d(9�6�U�f���>Z�f�"�|@�
f2�ρ����@�39��
��+����������J�X�}4�ٌ[�X6��Eh���˹x�q�ӎ����qb����.A6�z��=�龚W�P�3��W�;���Tˑ.���@eІ����L�N*�[��6��(��������b�g_�3�ޘ]n�֖���B�`�qE�{�.Dه���L��2(�c��p�%6D��
�@!V8��>j׮�	I�
��(�,�_R?�Ȃ�X}�O��pZ#9��]SC.�am���3��$i=j�zIϸ����7����s;����2�����Gu�{�?,ُY�khi�_��K���+w~s
��a��2.дc[,{���	��$X��C$�x5S"R�{b�Aٓ���~���q�?��+�]8������n�����B}y-�@-��Qxv�OW��꘻�f,̓D�]��j\E�O�	N�M�~����x6A?�q�.QL������%�ٓ�^�q�u���5�(�(��;6�i�m@�K@�?���lދ�S�/<�6,��z[|-75���e��h�Q]E����L~�Yva�u�^����D��V�;�'���-�P��p�U�A8.W|��&�ګ�����9�1���|�LQ��M�+q�pk:ޙ�����/�������J����wR��)�R�X`W=�>��=Ly_K�����("lac��I��(�ꏣJ{��ھi+SO�t7��^cc-�Fg��@D���Q'E��¢&{��\���_�YޤXw��3���bt�r�ZB�1N�\z�CkRe���������O�dpK6��]�o��~E;
���{��W�>�P�Ph엡�/�ՠ�?D�K�\���?�J��/N�nѮm�0��xW�����ƙa��T|����GaC@�f��ϛƧKȐP��Cs��GII+�{��\LW`�gT��Z=�k���ay��a��RL�U���Ƞ0�XӪkl��d+�)��(�SDKX�8Y��D�@=ў�v��f�r��DA����P}q-����2�i�
e9,��BK���V��y�{�s�8����CB�g�?q��P����w�F��+]��
t��ͻ(]���{�2K@�Bu�)82J⠊�RES� �HB�����ζ��ޕ�0��_�~NT��.'z��b��u�}v����#��ƉP�,�4�}/�YNr����7�ɗ�(ー�0��e W�k�x��+ئPf	�����\��ϵJ��3U����9i#C�h�zҚ��VTGT�+g`R�ף�L#��v��J�}k.B'z�⃱$%wr�6lګ�;𫷵"��[�mҷd���d��B4*�?b
�����Bz2`��*���C����+]�N׊�ܨcd}�5G\dو��8�3TQ���"����{Ѡ��䮍�ɧ�à��@�@�Cl��*�ih]slk1�[[AxǞ󑰮��i%��P4�L�]�柳-�Պ쎫n+%.]��'��0�P��	��y;G��<�]y����[E�>C4K�/&�q����GY�?NL���Hf�4" �i	w��ڭ}rg�J�6�5��e�̴Z4�ǵ�ݚ�� �<[|��ӠiJK5�a��_or�u(���Q`	� gI�g0"��8�y����S���o����6�A�>$���xW"��/�ľ�6v��QBX�Me�e��x�B��H�;4ɨ?�=^��eh�e�^�=�1�DK�?��H�0.m,��=7��~�"Q�r��c����@
<�`�{d¼Ó���/$����/`2�V:����2�͌�9��7�� ݆�K���/��P�`������m�#f��k�H2U�4����I��@�I���l���&�ϓ4-O'zL#� o���Y�~��M�kW=���w��㓫��ɅS
WmKv��Rag���|�R��%S��ĭNz��D�ܸ�]щ3&�|���\9Ϛ@:�%/�﵈g��? v�Fx���jTz���x�r����6�X����h��SZ��x� ҩ9b���j�:�v�������������!�T��ݝZ#���"d�b��Zl`D���J���^���fk=	j��V~��t����X��,᪟m1`���J�m90�E�7eO� �������B��V"t,�!�p3��p���L#:�\�������ֆ�|�;5r�����y&
5�`S�%o�p���3��ۭhm
y���J$P�PM&|Rpd�ه�/w}H��Ȏb=99�`Հ�*���}�ʯ�~n�܋���|�Q�T'>��Zt���O�ݘ
���ha�������A� �ӥ�(-��<S}�~��`t�����eu���u�_��
]'�B�O�.��C$�g|Ƅ��㄂�*ƾ{H�����/�����hNt]
�i~��:ŋ��c@���������|p�X*����F�>z�ہz�)d�����C�����ؙ�١��z�!�����t��� @!7�u�h8`u���M=ήG�ZR���0eII�{O����57������3+q����y2��l�f���u�"��<�I�h�T	�TN=�\�^!�"��N�I/�JYD� �*YI�U�k�88�/(�I��Xw�����/��bÂ^�d�-�+ =�ދ���Ih�Cr@�TT�.I�3��]��.)�oʶ�Z��W� �4U�*��TB=j���m��%~K7���d�+�	Օ��c@�鷗)�s.�x�׸�����>�
Q�G�0l����	IZ�3���
�k�qxl�m�'���/9	�4���ɶ�`��m@g�]�.'户h�p777�
����[M&N�ۥ�V�~pG���m�P� �D5g!1C��D���w����0���Ϡ�^�@��66��+��+�P�u;��2�ag�(56\u��Z.8�4��$%�B�n�l�m�%�^+}۔���#�tip8C���~?T�t'�x��Q��jM���L-Ǡ뱓�	�Et�X�ws�g4��&�,l�����]���t���3_�Z�K~����̑\9�Ĺ+�\.�<h�A��^  ��R @�%�#bq�f=���"=-��b$��*�����&|M�՜�ݺ�Su��$AP���VT_�s�t�"��毺��oJ�ŢS!n�nQ>{4�z�]�>�qqq��Ė<JБ�L�R��\Wl�A�+�kHR�M�ى�w����&_�WwT��j5�:��o�]b�>��z
���>�2κ����[#��@S1��������y�GU�i2�	��@/vk5^s�ؖz�w��%�<��&ty���sqœ5iG|~6w$�˄-��`�
�.�Q����:���'�6����4�=�Z�=����*΢�˶��(�1c�D[��m*�k���
�tDw�|�V@��M����fw.���9{1B~p6OT�E
�Ov��J����BΚ�M�d��.Pv:'-&�1��mO���G����D}���G!Q&'ɗ&;�Z���C>0O�Vg�{We���� A.�~�5�0}�6*��<��[_�dg�f��
���z�~���n�D�@���Tl�*5�Ə��R���ױL��S���Am,yhÄo*�i����Ky��#<���wO-H�L��cH�`�N�&]��+��UODVja7F1CX��������!d@�`�d���i�y�����?m�S��ƿ��*}T�&[$�k�@־�m'���F�9��~�}'�