��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]�����j�ЁVL �t~�����Ev��֖�	�
�4aV����D%8���z�CK#�R�Ą��z����vϞ�s$ؑ�0b7�O*��&Y��Mj.R��r+�A,��b1n�c�����
1I	h�oW�F�:�fK���^�ΰ�ڑUYTK�ur����(9�3��J�$����f�����Q[6�¾x��tѐ����0$%C�:Ȯ���m��d"�����4��-H��th��p:���Nc>lj)%�a���J�=Y�oR_Y�3�BtV��|�̫����u��jd�n�]�ʕ
q"9���F�b���{�!�!
�ț�@g�x��{V.k�S��M^M��8o�<Β���F^��d|\��Ǒ΋�0$h��T|d���rk��j�Mq����o�����|�B��"�h�R�L�ytko�C)w��8����{\0�����h;����X�!��
R�0X;n��!�'2��=��) ��SVǅK�	۸�[>�Z>�<���r4���Z�2+M��}1����$M�뜘�R\��������xA�K �;��ѹ뾅��
���˾�����(4����&�4~2]1�J��w�����8	9Ƨ
T�t|#5��:��O���G�Xb�0�s�������ZWL�ґ�u���l�]s�;���yl.~������(	ɔk��7�r��tV���U��|�DQ}�1у��WP�:N�[=L_J��X%m��,;
8���ɘ�
��(1�$Qm��o�6�0f�wԔ��9B�?")53h�/���*Ϧ�_��v���z+o!K���K�ْK�{���q�-�$�d4�O�%�
���w'����[����	��ݞ�vM%y(��#�**����;oO�K�2��`��@�^.�0�^�{�4�����
�����d�k���j�>��p3�눧��4�_^��p%k�U��ߤ�(9y�"lpr��2�x�\�\ʇ�9�A�2�.ƨ��Y�'�:�s�*�S͔�!WpP�Yn�a�i��`�C��K=6����U�� �ظ���n�����dKA#�o�db��3�*|�@_�n�}��o���67��
m�����s]E�cF:P���"kTȥ���7��$�=s�"2���ڮq�Y"<SO���E͙�����g���y�}�P|D�CK>,��uz��(�uf9�Jvr��#ng!����cШ��4t]`�hŎ�[R�Ą
,������������L���!R��W}��
���ؕP'�E�<
�D�'�P�X�J©@L���y����9yf�i��e�_h�.�Y,�I�� {6�b�������6�ҬZ���^��Z�+���՟,���B��oJ�����U��7R:@0	�-?� �9bҝ��:�<{�1s���$�)��Ţ����6���^B~����h���BE�GLg�|w�D4�X(�͡*S�5��a�kў4�S1���ּ��fj�E�����U@Zċ]���%�|	�z��K�sW�ۋ��>�~D�ě����a͘���Y��^��)|��ч�E`w�K��W��7/lV�Y^9`��P�/#�����o�0���>s�V�I��+��{=h�;�$�ǌ��]t����E�ə$���IJ�L�D6��r#C9�:���~�y�or�����+�Ϥ�JN���h%�Y�v%J��kXrK��}�]�?C�jJ�3`7�\��|����l�ﳧ�3�~+���d��[�q�X��c�(o0�P�eR��2�%a��.a�G:�np8�<�����NOR���G��E��@�(�)c���~�Z����!��Z�v�t��]������y+Į{\�;E,��V&)��v"�.����[�GGN 1�.�\1O�H��$���䟊<��@�f츞6ph���֝}*9�fxT|�0PM(
ZL�M#� Q]�����3��cQ&� ENk�Uҍ�)~\�� �	ȕ��Bi�����p<�E�b���ᇒ��n�i�$�&*�I�T/Qj
�P��@T6�OOKpg#��LBL�pn#�4�'^�8���mti��Ia�&0�y��i�8�8��q��kt��	T���T����'J��Ͳ�T�'�:@�� %�j����@l���)�-�\O��9_D���~��x�P"d�3�^�&��`Vɽxa"V�:(d���	QJ�fP��Y�ҼK�&(̽���:l�Q����V7��(d�Sv鹲�Pnq�����AH|�$}	^�׶��@J�����d,���]ϖ,HK�����Vk��.s'�8�O0	�.QkQ6#'}U�����ǭv�F�AĆ��Y��EA3�L@R�&�Urw�j<��n^ #�Z*Qu�^��p�lR�U�M��Y�Ba~���Tfg�O�nzS�Òj�s�l���:��Ӓ��l1htM�obT�\l��ȭ�yR�7����Q�����U��}��)Ӓ�����^�[TE��
�������^����� ^���/�0��AX�>2���Q�c����>ϐtqRB����IKX#��,���D�iGB�+����
cA��5-I�!�_vJ�UpQ�/�����2�%�#������??����虪CX�Q�ό������i���9�B7��7)^���^��Q���K�����B쥎����5�]�ېv�t�R	i��ZCG�t�7�� �a'�����rq���F�N�)��.聙��w�ls#�:�L+���p:�Q����Uڕ_ת�(uF�~��5Pސ-��&N^�S²m�˾��h���NR��5v�e�����(���.� Hb,qЦ�o�^&�s&�7� \�2҉��R%��ɏb���t܉�t��h� oqƨ@�3=ߥ��)�p�������ƹ'^���in?b�Z��Y�Du����*��ܻ�|*\	.�$��2	xQ�'F�E���N?EH�������Q���VA#�MYг��(��l���/.�����[�7�H��*y4�j4�i��+����&h;�9�R����"���J���u�z.�:M� �����r�-2Z��{2!l�Cnn����e"��Y�t[�O&;S�.���O���Om?���Z�١)0=�j%�M�?3��	B�n6��[R�����|�v%�mA�S��Ѱn�%��q�,�ݟseSj^R�4`�2Y�w�Wbd�$ ���ˣw4d����h۱���)B�����7��~����ϥ��P����#�R�W�j��rf-b��s��x0���I`�^�\��qv�!��7{u�E�|�ǵ� ���H�[8� 8�E3d�Z��Z�1�´�鹎k*e6{|�����N7��DOJ�	�m	G;�Ӱ͎a���x%��Z�w7r��X�$�T$����|<3��F1M�s�yD�Wn�������m����a�e��z�g��
�'�cp��&P8�pp<�L�W�tر��p]e���?�AH{�b��lc.��Vq��ml�ua�yT[����W����5!Ė	� o��I[|�;�8�ca�y�橊6O�����'�U���av�9���zÂ�ȅH��^s��v�G�>���X��i�ot9�N�j�B�9��8Jyt�Ir����49�{ B�/[ ^�ݨ�ɵ�CV��]H�bMu�VF�;5�<M8E-P��s�u�ɪ���H�Xy���K����6S?n����(24�#��l�l���M�l��>��z[.`E��?.`�N|�S w\��ͻj }�}g��Ci؈�Ŵ�W�Ć�}̐��M��XK�V�m�U�3J4���4`!�t����'4��esU1KJ8����`V���R���d�_�	$�Gݴ�N��!�مtzYWM�>���e5�=���_g�dι�U��*m,P�n�X5*ZLs���ȴ�{}&\�ь@�MT��I��}��>!Lez�z�|K@Ӵ.6����^L��!�腰RA��=x����r��H��`�k�X�p�)E�xR}���{#۶Sv�~����뾙�L��Db�ݹ�̻H��8X��ͲM���Ae?�ȭ�/$`����Ώ�p�l��*׊7#�z�&&������W�˅=ʑ��B�5;nҖ��Z��r �qxb1l��~�zfA�,�S+�MmS��d��j���Au�4�T�B��Q��c����4uy�_���_�P�jɃ,��z��5��2�GV��[W�71�a��#GaP��x��_�(K��GР��c���W9e���Κ#��j�����;g\�����j��̫ϫ6E<�3�'��yʊ�����Vm[P�H�)~�Ya�D��94��X�&��C����o�ٴ:V�Ϩw�Oox!K��΂2h90]�#��J�_Tu�`k~��a*)���P�O7�\��l�,X�j��荟J������+���p�Dw-�E���V��F�w���䠴�V��Ă��Y�D�gG
��]>�a����|Xd��x ���$!k��#���K�t&p#�a���]���Ӻ�Q��V���������N���y�>�7���r���m�u�rz`>�x ���Ϋ�2I��5�hB���7}��[v�������"�8ʋ���������]!Ӵ���H�_��b(xR�Fr�]�0mwb��h��nl1d�=;�?8��T�����/�E��'P`���e���lV�Rb�C���}�c��B@"Ǫ�a(8�6״�F�,�`�&
昳�S�^��^�8n��ʹ�����Lod��r1,�eD�=ʡKl5Bη�⸳3�������.9j����N:<ſ2k���]|�!؆��	4KS�T&�?Ų*�)�I����
8F]9�Wx�B-��O��D�Z]�@(j.*��e
Ԉ��R���V��q���ꈆۼ`�>�ļ�d}{���l.�UKvP7�x9� ���o8�D׽�,���z�5&����'l�iH}��xT&?m ��lf��ξg�c(����&����q��.��b!た�Q)1��{�4ɕ[�1��{��b"y�tW),�|�u���G�?>n�3�:j�x�p���tȚ��i�r�\��>�}$�w��T�T�::, 22���#�u���GZ�+�40n��m�s �
�Q$���KMپ����j��Z*��E���<� '��D�+jʅ]���L1µ�e�Q��O�.%&K*����m��+�7�S�+���&C>�<֒�O�`=����V�7e ��6yB/;�B���/��`}0x�����Q��5�x<f~�|��i� s���7>�(٥=w�qN��������G�`�ִ�NM��ՕlK�ԲB�����3Zȁ`�O-�9���)ߌv	�P~�5H~;�ۯՄ5|�&���ϰ����pӊ �mu/X�j�4>G�j���a�К�t����C3H�`��G��^�B�#�H�y�L��	�E����r<WY�3��-��-�zK��$�ֹ��ꢣ��b,�KڹP��~�.�u�x�ZN�U�OG8�	��˫R����WL���c���Z�=�O�q����:�}�OT���׶[�ȉ�:|�sj��T�.���".�F^�\򆳵��0.�B�@i�{ �7�����PoDI��^t}Vr��5 �"y��4��nK"���I��x=]>���Ŀ%j��$k5���kr!
t�"6�Mk����b��|�3���ݫ�S���N� ��1��wE�� c���ԟ��=���(��њG,&ԏ�����XR�Y�°�ޥ=�?M�Wy�4�x=��Y%����#��4���~7��Z�� =�x�7�|a��/���q�W�p1����js���-�mne�;b,��j�8���"w����v��>�^���L@��GF�|ؒ�De`�b�{��d"��� ��]�ŷ���4�W�S��C5i����(�dO~T�3+)���5�+�PaE�Fq�9�R�� :���t�x<�eTϰ��eMy�^�dR�5p�U�d���B��U�>\�<�Y�y�ʃ��o@V�-�MXz��޿�&�c�p *�{�FP���k�~W$K�"k��"u�+"i�s�
���X��@;*Զ��m ,ŐV.�s,�\�_�m-�X�N�H��h�ɲp�?Վ!��S�<�٣N+�uÄ,�o��'
"V���We��ăy�d� !.��:u��Z�{�ݮ�sF}ηb�&<�>u�������n$H���%���:C�$�����t�z��)��ͬL�P�4;������C���_�~��P�f�p�5g�r��I���ѹ�&�O}]�J=wh��|�d�AL�� �
��[��ޕ [Q5���|п��x��t�END/bZa�3��7���"��׃0z+��Ծs�:�-PH�/�!pk���Zl�qMb��X��a@&P��x���_�y|�kP�|��j4D��+�qp�QЕ]<���Ok#c�r[�]x�tXt��VhmC�����a�	�\ ���_�j�+�\�5-{��-��+j��vO����V�)O����_э��n1�����pӳ��
�3��ZLw����`�T^�"�����FD�ZG�o���\��[8E�Q�FJ�� �wu��+�y5�ԫ򞒍��:x;�}�yA���]C?b�.�&;�b�:��1�M����~.��%x�0o#����'�^v��i@�d�׫'��~a��?��ͻp��;U}8�W���GHq䀳�;6�5O�ׯ�,wЎ>w�Zn!��V����a��tغ�x�;��u�D�OI��2�h��F4�W��,Yg���t�g�N/(�^q��n�3�1��-��bV�`�}Ʒt�|K��i#m�Ч�˿���&��:܆�&�#4fw���@��M��c�	���xr71��uHK�_1=#xџ��ܷA�������Vcf�@#�m:�:V*�beC�,�V|ϛ�'C��v�;ݢ���	U��Q���n"d�l��#�F��,W�wN��,�V�%;a�����Dn�%�!�������'��D������]5?��,��a��)xŞ%��[�H��Nez+�K̋�0���\Q���� $�
π�9O�j$e��#�ՙ����Z���YIS�������.J\0潸����^=�����D!��ѵ�zp�uC�x�ۧ����Ԛ��s��4���V9K��d/Ү*]�*SAD�
���-�[K�p����Ɋ���A=�#_m�O�^��8�د(/eԢoH�
}}�ж�ĝ����<#�Ŋ��{��O5��.n�~ ?�^����oN���,�	���QT>x�҆7V\I�<4���H��R
���B���S��] ���T%H45��h�>��c����M��KuI�^�7����jXW�/���H]@c��	�W&oF���|TB��@���$�]����'ޗ��U"�y����e��}�E�R�eF5�^c��`|����S���`p��f_�:zxY�<
��c"�P��
��6=�Ic<�;��?,yO[v��i��'�չ�;�y�M�E
g
Ķ/2��Ll
�C>��d|����kU_{Ț�E/Ǌ�o��=S�2�Se�������.<�V0�Àj:�<][�!x�}(A:�}�Dއx��w��MK��v49w��'�)��K�>Y� ��h09�Z+�F�F�_	�[E2~�:�H����qd�����Ia*�g���C�16x�3D������:�#��} ������B�Ç�aM]�UlN�$bB��ǡw�*�����5݌��=i�W�#�&l��pU���;ԡ=��V��+�-�_�$���
ݡA�$�ꈅ&��Y;�;���B���_x�Or�T�vY�-��PUvT	
�Ϲ���ӤM��L�>�N*���\�N�բt#|��2Z<�j3�{��l�����~�TC��65��?2�{z��N�F�H:t����gG"_�[dC�$��Jχ�*R4(�#��a�5Ne;u�[�͵�*)�;���l!��5���8H´]�=�����Ҩ`�/m*�l}�'�
��!�@	G}�=f@aqIfD��֚��F%o��&�	i�!úF�][�b�XX��s��6�eNѧ�ͭ��}щ�-:K�3���L^�h�
�;}T�즆�F��յ-�k�8K7t�����g H�&�4e]�Q=��%�ZR��%��������N��K������ �AIi4Z��fnMu͜W]� E� ½��a$�P��􄂄#2/�W˭<�a��.Ի�9��}�u�iEʖ�����_�yu�e�^�H�/�Q���l8j�fEX����w��4N��!�h� �M:�{��O�m���D+l�(�*�7&�/��� wJ����N�ZT8O0��s�g4+!�a��5o�L�,'Z[�'�e���=k�:D鰤##H�16�v��H7�Q, �ՈMʘ?V�[z���]��1*�
b.T��/I9�������s��ko8vd�mұh�
��&���[�_�!n9�;Y��"�>_�Ą�yC�u��5B��f�L�VqZ4�t� #���t���8C��>�;���Ǫ?�H-~���Db5S��ܼР�c�D��&�S��B���b��Ñ!���s�J+6����Ryr�mnh��P^]^2��۬3��5_�����zع�9����,LY]_2�6Ù���s���}�`v�#��{�"kgi��AYr�h��R۠���k'�8k���zfq �b
;B�t�R_wɁz��+�S�,fa� ��4���*�PŰ������@f����C��ùo�s�xM�]A�PT�d��?��4{�}ԍ��ې�Q���E���u��An�!At��t�>�ò<��� j>�%��]�/�xj�+�ɭ k'�*������N_���./��uK�H@"l��5�Xp4�s���M�)�L�-���H�t���G�!�,{^�z��Ck7v�D$29~wkt@D���`�&�2#��+����u	�߳���{xF���|�+�[V�gYj���b� o\j�o�����8�i�ɋ�X���Փu�V�a��yz�Ȃ4$04�"���:e�7|C�z���$-P��{vQ?m�FHڢ��Z`Z��܍k湘S<�|X8��}�B> Kkh�;ρ_
��3��`O�J}�"�\����1%��qKd
Z;���5g��/��>J�骃���h{�e�O_/����7G�ߍ�y��#A=��M��S�敲UA���_D�	ʯ�%��7���'�e���f��([��վ%�Y�δ�i�Gn�IYn%��ȼi͍�@ᙳ6�7�SsU&��a��p�qU�MxD�ց�)!x7��[���-����_�YL����٬��ROp�	�v�9.`{��3~`h�`�J�n��D��*�\����]��&�����x��wV�t��`�+��P�X�&�h?s���ž,~�+�k3QJ�����~Il��5�=��Q.�D%��X���K�����xb1�S΁�5@��*ַ+�U��V�ʿ�������Y/y+E/��{��!�l�:?�T[�e?�<���eGB�y�0uV�c8�iq.db������Ā�N�5`�bܠ���I5!�6�F�;��;���H��c"2��6ڞ/(��1!�#HO�,��Y VV'>�?�ۓ��Q�	=k>�z�t�e�fF��~�$�ދ�:WZ�Ws�_���.P�z�9 �G��i������� �!*�W8���Z,���+767���[�ԑ���+A�'�	1n�d,8�.�'��H�ege/�ʁw�v�=� �(��,������>��k�!���	���s2��xl�b3�K{��+~a,⃕�����oW��j�Q��5�<)OSAt�8i��: ��e���'?O����7Tv����t�BW��}l�,,��A;N?�T�!,��^q1^��C�|���8�֪l }��)�j��[B��>J�����&y������Tc�h _F<�D�=���w�Pw67��e1\�ZA�V��\yq)�0hdZq�M��{�Nr҈�f�����m���w���肉��^	.�Kk�����k�Y?BE:����H,�H��@�����_���4�c��� �S	@әv�#������&�p����'�lf��;�"���y�C"N��E���Z��� ��f�v���dZ?D���r��P���/�آ\�"dܥ�h
5 ��z���-��$�Au{��9�)���Y�������P[�I���W���q��-��j���-=i����=�?U4>PH*K�����7�}�U�	��r��*v��T�"S%��j 9�����R�Rl��s|�X���d�iWC���h�q1MG���r���h+g>��Q��H U�����b�s�_�l�t�+x ��q��A�"�e�/�ݗ)��8�y�$VF�թ�	�x@}i*�e��g���`�T����-Jb�X�� |��� �@�ß�g�<�@/��\�HkJ2���Ʃ��ElEZ������D�.
n '¬��]���\Rq�!� v�j�z���[�`y.�I0��˳f��9$�2C�
�`�Z�ؠ�;�7΃�Ԣ���,�=O5�hZ;P���SiK�,�lJ��rIcld D=�)�0�?`j7F�!mm���۠BK�~	+n�=�x��q_L����k�F���ӕX��Te/ܰ|�wq�ވ�f(Ѣ%�9�3�R���I��D�]@���\���3��iLN�B��=͝�c�������]��/]������V�>�BDɑ(z���#q��B:[�L���8b`L�31�_�^<y�}<xg�"-dG��ѷ����o%[�'Wc�16~��XٻTp/�v�C���� �[Z�����ɐA�� pϦ���k�,qD�Σ	3�����M���Z�k���O�3jz�?���v�A⤊\��'c����J���OE�sJ���Z>&����E%� 1��}1	�eĘ�T����xj����0�[��:e-ͻW� ���(mJլ�OC��lc`�����p�� ��yy��''��w�����&�ފ���K	U�4���c�+�ߪ6�$��|�	�>޲�H5��<��9�b�%�}�qpZ���`oH�^��Wſn����t�B���/^�V`Ѧ���/9N � ��CF�Q��U��o������ݗٴ�)w�B�J�)F�LYs��a�PL�ĭ"�	R��5?����c�������U����" N<PFp �YF���CZ�N/<�ž`���֪-��V:D�
1���	*��	<[�auCr�Q���Ɠ�j�v��ѣ���¥�e���M�
������c�����ZD���OT@�"��m��U_�f,`S�#�9�5 n׋ޠ3Ӷw�޳�I?��P��d5Xbp0����������Y%iS��V�yϭ�5�=��D��o�uSm�`�
(���O9��k0Ƙ��\L$���ԅ{��2&�d[�{��������Z��[��	���Y��'p���Ք�I�L'&�����#9��1���w��~C�a��x�����������_n�>�:�az/o+�n�#�<����Bf�C�5$�� `�*b�����)	�5��i�m`ӛ���<Q���H#mv�r�s�M(q$����b#�3�7#�5O;".�5,���G}) ʘ��?���|�0���2��6�7(n����)6�ְ��忇��ƺ;�^���N�^D���]<�	pm=�c���M��8^�TW��5�����&����P���,�%��o���L]'�M崸���L�B^�?�,��T�e���Y2"�:�rty�)�g������%T䜙��L��nW�����]��Җ�A����u�)����G����<Q���᫅{6�ٸPp]���k�S[�N���y��6C���T�I|g�QZ;���	_�+��B+�_[a|�)���.�	u��t�P h�<��+��h����E����԰�5�O ��iSrz*��nN�Ĳv񾝭8Gی&G`L駟��4��!��aXIdT#�\l�p�� 1��@���ҿ.�I�p�a�뵚�C�.#�u~�8�^���	Z]=̼��"��,&��ǜ�(i>�W�0�h� |V3ѴX���Ѹ��sYľ\0���>�9+� �t���Tghں�W�<���a��jʑ.rW?��p�j�蟳���X!;a�/�����K��n��寍� 1�c���=<���-R+�S�_+��ly�q��VX��8�.4��� �k>@�N�����e��v��eT��5	�,�f�]�A�b���y?����OC�>p�S��gm���X��ϙ b��FtzŒʆ����C�Q�z�r`E�2N�A����X	���	�t>JI�^�ɵ@H纟='�@�EY�u�{��U��1^j�oO�"f��i���-þ�&eӔ~K���>�ϣ�