��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����Y_��F��tw�p�^�=�����DW!of�.��"�"V�8��Ua}W#R�M�-Q�xq��ų�����#k_Q��?���B8I��c��l��{ͪNȽ�D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����~�Yp����ƅ��*B_.� v���z�S�����đ�d\7~��}j�T��z$w�K�<�7�P�i3���@����崡�sU��,��aN��s��%{��u]P@�~�2��e�@x��=fG�8�&�F��^��d�(g�`廣0$V[C� ��,�&�A�t�ə�	U�2���\��,I�e��ׁ��ѳ6�d�b3�R�������B� �ć�&�40�6��?W}�B���3-3����XC�����5�T��7��6��yE3ӗ�p�?{���r�hu�3ߣ�y�X�0��[�L*j��n�7���h�8�F�����i�/��S����*�5�M9�=�4�P1�S�g~�4�L����W�"����۞����'�4����Bl��.-�SX҃):gۈ���aJ7�st�f�r��"���Q��?LGs��Z�&{���z��G��.h2���%���PU�O���Xu/SL.��QJ"��Xu�MYW��rK���u�v���_�	�}>��f�5C�;Tmr�~%�J:/gQ��,%x�3%�޴�	w�8�8Gy�Y*�#�<�d�3t㡥!x
��!ք>n~�޵r�m ���##}ö���9��|B ����H�O��ҭ��l�8����Y���:�)c�<_a�p���>��z4��1=�W�?����*O���X�cH��r�j<��8��h���P2�(�(�c�pD� NE�e]�˰?�]� I!�>#��0�a�D^�r�a�.��-���*�^��m�Aͨ=��I[f��'U�爼��+������(��� c������^��g����)]����ڑ���(q㭫�4�@��$*��g1��F�[r7ϧ��SDS%�ӯkq�1A{�1!����rBX���^��-r�MZ���ꘋ�#�M͢�o¼H�����P�=�l^��"(��S!����\Aȡ�#�*���쇋x����ŗ���1�A��rrU�|�&�����(����V��MsW�	I�����خxbyW.��"Xi���Q���M���>�[s��+����JU�"U���Hb�����	4�m�W^Bm�\K�*�h�Ga�r��<�h[��rg�ʚ����ψJȶ��hh'kY�]�
)c��!��|�߰h�e���8X��#�-���W`qf�7���氦z�������=�4��:mFL��;�� c,���Vi:s��6��T�A˨uF�W�5����
m������2��Sl����W��w}��y�H�����Em��%�\�؈�|�U:��R_]}�ނg�Dx]���&c��p��+�Sn�S�#�e�����B�Vv�[�vC,���SU��HQ�&{���V�yP������#Kh���\�ߤ:�������1�vy��S��y�p\eA�d�.�o8��y� x�z!*�Bt��/N�����W����q�� Э��� ���n�p↸���#���T���I�@e�Y}�,
	����׋���9P�u���[�W��D� fl~Ǟ�T�P@]�d�L��P K�F4��̍�w�s��3_K����s�-����[��`�m
��7$���cؾ8���ϼ>���z��o���`�~	�Եɧ�8�
x�K�C��(���W� U�L��n�"��+͠d����:������Y��{zl���f���2&�{�j@��svu@�@�����Ӊ]���\�2���p�~����`��2ڝ@��_���S6}�����G�'�B����ȯ��6&5U|�H�C݀���V�:��bń;�fc*��gK{�#����(l(NA��P�_�t����$�������sI`]����`�W;�PH��
��$h��`��/�a���)��E&�v-É��� 	Z-d�M|^9�Rr�9����s�=Yn���w�B�����N����pX��֖6!\7������ۭ~�B׳�$�o�d����I)���`e����y���Vy|rR�e�K�_��a��k[m�����GxB8rJu�-if����K��!��)ی�B��(&�D�;=;
Eu����;a'N48�Nht�-����G���W
��rfa�+�o�K�Y�>�����Bd�yy�����	����dr)٪��+���r�c��<D�b=���I�_C��x��l�h�>���V�ݰ�r���}�i� L� פ:]di�f��v�v���/�X�(�F?�3� �S�����4.���ϖx7P@���Q��|4�c�6.���*�����m�8
(yX+�:O�q��
(��gȥ0�[!��B�5�����  �< ��|�|���s�l�'ak�tz*}������)E��$x��O�i�<������P�I,��׌$oC�B�aί��:���U�$8.̈́�����0�[Üsz?���ː�_D��ch���؜���Q~�'�{�}}�1�>^�Z���Nl�#�i��4��w����J�EP�P��E�ڄ���{���H�U���j9H=�M��F<����Ӱ��]&xU���4����vxG"�]�m�P��f*���)��62�E�����l`��=�W1�p����f��,�!����;�^n!iiG�������y���4�V��b�`���Y�b���O;5F��h�R��\}���M����M��t�]aP��s��f��&א��3�kc��@S�燇�N璥�������ׄq��ƃ�UzX�^#˟(Y�k�<�)E����;��=��ך0Z}L$� '���f#4�}6�M�O[v?����`����Lm��qop�<ȏ��_���X�����`���s��0���G@z�0A%,���U�[xI��[�&��E��-��l��.�3%�uu��Dӻ�/�n���>j�;��o�h�Y��~ )S��|���(aj�.8�宄��˄|�c��X9�O��S�d��$ N��<�YX�ݞ�¤�;�~,��GҪ��PIo	���)H�F\v���N�i��\	=��'e�_�a��K���ްY�$G[�],�z"�>�"wE��mһ��j���U�R��Q�]��&�2.a������Wp�IvX��ֽK�p:шX�j��z󴴙#�Lp�oT�k����p���e��Ұv^U�������G����tj���o_�!X����|s*|�b�$6q��:+!(#뚠b�Z�S��_�� �uP1�ދb8 �M)�I��JYԧ@@�H"(���d����"4��=%����<^��"Z�}�w2���2�6��Q�_^>�)��w����s�q��5��ȃ?�a@�f��v��^*�YW���]t����O 鲬w=$ٖj��,�5Yf,7�Nf!�EM�%�~�h��4�~6�R��t����P��$��!��l�f�i�Uo��.�X�Zz�R�aԝ&O������(�ې�(��X �vD�@q��_]3�<8q&Qm��Œc�J�8�17�2;�^AD5;/o{o�Kճ.���b����~~����u=fޝw|��-�ѳrY�%��=f��pR�l�cN�ʽ��ǜk�n���Tm/�����$0��K������W�'�}3TK�_��6�ێ%����m̼�iӫ Hb.t�e<t��f$y :�xċ�b9T�L;-��^`�ao����,�O�CM_h�̤F�􏭝�s�a���`��"9��ҭ�~��z��!u���d�x��hw�=��~B��䳈�+���I}g4������������\U�����Yc �M�4���
�ˀ'U���:_8��4x��X��lH/+�d���D���&�;��㋹� 9!~�1�Y�8��b���EMU;VԢ�	�I϶[���M/4Z]��iX{�(�}�Ii
Ez���py�eО�YubX};p�@.,��^n���|�i0T��ǅ�	R�K����Ep˝�#I0XőO�W���3��O�wd\�������8������
o#��xߵ�s���i;��Rc�v��?#�e��X�"?>S�Rz�/q�,����$ ��b� h�\/),Q=�I�-�V)g����`$��ѯD\�t���Q�"�<�����9+���F���!���$hl�U~c��"�@�T�Y.���������{���*	��Z6AF����\3��0ş�A�:��Ƨ��"�b�W�ل�c�����{4ɻ�0��D��
2�9�}:���z��"T�f�%�BI���Q��R߫�AI�0���y����h5Օ���|/Q�v�8%wr��5�@�����{�13����3_�Г,�<��wa�#��%��.��y�����e4x���B����>�b 3�kf�����x�?q3�f�����U6�=�Ж�I�8��BAM��`�9��_��������RYB�jv�{#�5ob{��P2Y��J�.�j��¼X+|��gTJ��u��+U]Ÿ��ʷ���`�����Q����-Aǫ@&�%�OQ.N��Ӹ�3:Ъ.��dd�1�fЊ
)獞M
C )��Xl׉��&��Ƀ;�����'�ivh��Ogd���*I�ʂ_g��D�{����V;ۻcX=��֬��p��
��-N�����J��"st�i��W���մF�����hw5� �S�j[q����WC�_/�iO#���:��I�#;�1�WAv�P�4J���$�3��FU��f�?ꙏ�L�z?'�b{�q�k��7��YAmn��2����RO!�_TP�!��FO9�j�~	¸�&8Ov��mi�
�@�B��U����2�ʹ �{��`�X|L�]Ċ��uI%k+W |����%�1�S`1t��r!k�6�8��U���L/0��e� ��pW^�4��c	l��$��H��'����[���*�ӳ�r{g�,D�'�K��'�{�NA""ޞ�}{� ��Rz�r�T|Q��:���s�!�3$.�{��MO��X.W^3�F����@�1�V��k��M��#�z{t����҃0�7 
��y�v�4�	ZB���Y��4�D����͉h[�%�%*g�B�Z4���6@�3Ð㐗��M�^ra?��%Pi�yG�.�ꞲXj�b��1��z�a�N��[�ɓ����̠��,��M�8��E�u�{R�1�Zyy���|�$�R���ԩ.���j� �;����֛W��<ƭ��r�����!�`{j�	@�x�(}'	����#	��}^姦"��F�3�jQ\^`H�W��'��Z߹(���L�u��Y�j�6CD�􀘡����/,�zHxL��[P����LE���]����x��{�%\+�DS�*��Hp#hT�EW �6�F�]�H��U0�߶.F�-R�w�69��ɜA��u�.G.���*fSB8����aq���k�]�iZJ���o9��d�eG�u�*�n|�|����?��6[j���o�_+���՜��yߎS;�Dm�KȐ�5�F�MLt�B��H��u`q|��"8d���B��q�Ո�Y#������\�*c�Z������ ��CW9�!m�JfxO	Cy�h�'�HU6Q ���mh�y�wӥ����F�����F����A`�S���7�5�=%
���㹟rL�;K��pJ%YL�֢���%����l.׈F���8�,���w�oV0���j2�Y(��ܑ����P�rr<�WA��ɫ����o��(;݄�Ax�ĳl�3�9R�1����R�27�Kɖ
����3��ɬ9>��u�۵J�}�,�I�NҸ�b�E뭕s���V�Bi2 l5������Y�["&�%,�hqqGʻ~�T��U�Z���j�PJ����Ĕ}F��:��8V�;�>Q|��O�3[��M/h��&��6�DF��L��핧���Y��UV�ǡZt�ɺ9D�ָX�Z��~UT�Ш%��ۇk��.�F�E�ћ
]��d�@����e����(;�oaն��9����!�0Ď2]ta��MGKŢH����|S�����mso:����e��W��1��w}P�Dr�P�U��ff����$��y���y?���&�d��Qշ�`���������~�υ�2�T���i]����c+�8���H�U�.��I�'^	t�C��â��0��P�a��t�Q�C��_Ep���d;�(U@�s�ʌ(|%�d�$�~���{\9;[V�C�c�f��#����{(\�\�־�Ʋ���i{�!j ��-��P���X�a�΄������.;� �� '�$z��e��m)����֫%V�P��V�ܰN��hx��ʻ�<U�
�[�y���;�#ػPx��<�;�	v�k���4�*��&ý4�е�S0w і���4h���Xw6t�_[-��*Y3��]�YBw�ӧ�y�C�<K񈔖����Vp���}1����K�0�������7dt��Vi6�� 1���� K������k@�-EM!�(�<pX��]��=!U*�:��5��C팹\nR�OJ��o3%$�L;�վ] 6�0U�d���o��I��q��^��B94Q\ �MXp���ZQw���]�H����8��X���b6��@DG_#�N�Q��;�Q%U��{X!9>��mB���[ëO?%H���S-��@�\;�Q��\���%�8� bP�ܪ��j,TlY��7�����e��1��D$�͉=�D�e�����&e:Z�`��#�
��D�f�;j��l����K��a�}�mb�����J>�3퉆�Gj�����ӈU��������Dj[����@���!q���D١��ɴv�v�uI�7R�R����~������C�8ޞE������q�o��g?�4q&� �2��?���uV!!�;���E�����-����ÏSKX6�#�i,lj�c��3��j<&W�B6��~�k�es� a+�gQ��(��=�DU����a��_߅���]~/a<��!��p6
�<�ڱ�;�	��b)���dJ͋�x��(c�.�ܠ�L���˜�p{h0*g�y����E������Z�F��~3�@{�H���>���>��<�O�I��,_[�� �x���#eDwydB��Z�OK����Us��*�6���Ed5�߁���A���DF���p.W��A<q�i�Yp5V������?f���!�q�;�]��L����>S�"������#�Za�-�.��d�V��}$"�+N�Pd�9BXo�7YIT��Z[+�����Ӡc6q������V$���IJ��Z�g3�KJ%y+&�;a�>kExį�$o��<1u�K�g��z�������?%�qT α�{�\ �W��Y�u��_@��%^�]ߏ^�P�nέ
d��ʯ
���k�^`2;aYȽY8��XE�&�"�N��F�Ƙ�@��� U�h3��t�!t����2̴oUEg]�ii]����P��%m��)�\�C�Q�)�T|A�F�'վ'NT��Ǚ��݃�J��jO`Q�D ڦ1=�����N5��GJ�����ֆ�/���|�h�����zC�'�v<(����vP/�0w$�d�4)UGM��W��n59�lg�Y��auD�����c��w����@-zZ;X�=(u!���q����̭ZUi�BK5H��S6u8�s�F&SjW�B1��&��C�I���i%�I�2�E���M#����Û�Z��� � :ɢ�)Nb;^gF��#'���h��_ov�AŰ�����]N���s�tJͤ�4�dr#(��r�����s˒
6�(x��T���JJ����7��� �C�`6�a�MM蛷{�g�vd�xn�8�M{��a>`��,�
��:���5�e��wV��b��oq/����� ���,~7~g��M�0�3���b�a� g��\M�ǫ�m-�:G�Ԁ� �r��g�&��??+�ʾ�j�ܗ6�����?��&�R��OB?z�hSQ���Tyc!�lfs��`�G���]��*�ْ^ɢ&� V�����{w� �����[7)a�B�m���Ī9��[����7h�� �eJDD4_��\��le�-k<�P��v,�[���g)_!&�z̩����7�\��噄�R#|���L(�s�NL��}���u�U���F�o�a����,�٬�=r��%��3�$F\��p�I;�OA������h;���(
���$P����&��-L����nĂ9Z�
��.7�^�9<����ݡ�,n�
m������H����� ���Y㾪�Ko��c۟�|�~�>�t��5Y(�����:Q4��L,ݞ���֘�1rns�$�����c}�>��qs=�ȭ�Z����ڝ��W��kjtO=�ړ�!j�nee8�c^@oJQ�ǭ��
�����a��P�ߵs}�+x+�b5�M5�t$Ep&�J+�����W���׼/�Sg�Ym�֬�vg3%v ӫ��%��\Ƶ�ށr����n��P;�WD]�?�[x�S��_���P|��MWTp̔Y�����z��F{#܅+�B�륬�W#&dV�TV� #���F�Gi@A*������}h*��C�����e��D�ƚ4~Hi+�W�M!3ꦤ�4�����U��m�Z���,�k��(���#�"!>�� �@1w[�� ��d���!��������҂��!>��lXE������,/gL��� cSf�Xb��l��" CB�0/��)�҆7����!�!M�^�}�_��"��
1�4�N�R�ə[3��2aw���{���,q"uK`@� ���`-z�+��Z�� �ECN������R�M�|9����<���_p����t�RgEpd�e��n�I<
m�{���_İ�����2�F4� ]Gӧv�+vv)E-��(a�1&��A(��N2Y��R�t�9
YG��2AR��5}?�}!)�'hq��a�)
S#���Y���`�s�X�R��#����m�*�6�7�FИ���33Cޣ��+e�KA�\&{8�g�{8�nk�+^[MZ���ީ��Xj��1�v�iHdD$��F��)R�al��|���i�!M���MK���p�^�B�����<��=��6�*~��B���n���7� /i9*��
�"��C㘻��O�}��s�{��Ъ�<�U�D:ς(i#�Pic��$yv�ƨ�6Rw����F����ӎ�1f����r_|	�;������_�$e.�3�����^F�p�U�q�
��7�xFEv�!�,��^U'ǚ�I��6Z���3MX�y����έ�SԈ����������X}=$o����Ӫ�C	bB��zڻT�&S�f��GrHu��Ѷ� ��;����)q�×cV-�U�9h�w����s�8�?�@0��|A�w�t��΍$NLz
BwY�*G[�s{ו�˔���?ۘT����E@� �	�:�sI"]#wVe5e�)�U�M�-	y{zi_a�V��2ը�����xI�j��%��y뎮��-���r'[(��<��Y�/�*7zP�]���4����>Q�5�����0M^�vS5*e�,�]�*l� ����T��뒀̇�#��<����q	-��K?�TL���Z]I/WQNk�r�'� ��_cM�~��:[>��Ÿ[^:oKEH����SD�.�甠t�n���I�B�f�B�Ɇ�0�q8���͘
�r����?K�)p��~˄4'��{���ț}��'����oG��h��qW��6!�� E�?��) c7ż��+��&��z�l¹IZ��&D�>��H�&��̯2�h�����Ŗ��1�6�g�0#�U͈)��s�C�=;��a��O��?W!����J��OV=�]�ܡ?
Z��s�X"�(E��4�'Ҟ�����޴��O��b�UY�u��(r�ӊ�$�^ύd{ښp�^%�o�G]��l��E�
_|��v悇h�_��J&��I��O����'�ջ1Z�H,���p f�� ��{��ӕ�ḥuҿefL�������A��-��
�F��y��z(�|]ܡ�B���jهM���.1�ˇ��!�{Y����O�i�hR��.�ֈ�����
���Cb�|GC�ڗl��:$���4�)M���1~K�
#]S��V���Si�/G�BoC�h�%�F�_yR!8� v�ds{)��D?@O>ĳ�Y�=�6�U��^���8/Vb�.�����!�,G���'��7~��}�%=˟��������m����?�k�NK�7���(ʱ�ɣ��C��bX�%.��I���}5�Lπ;�v���la6�<���d'�d��6K�zPN��i��,��<�	��TNG\}��U������	�Ѥ���l�%����q-!����H�춾��=v�ё ZBT-��+����(�珖lY�Ƀ�ӱ�f3AU�	�^���B9Z�Mnx!j��8�>���qB�*_"e� lQ���<^��%�8sKV*s�k&��|�7,$�q8�1��Ƀ��P�qw��AQ��0�؉XHZ>F��K���
!{�.��P�H�I�V_拾Cʂc��k��3s1d�eI��>��J�D�➬E�;ӝ�,���s!�TЧ�pUl�d�-�$�Dt�Fxn0��>����t��6��LQ}�a�#�փ�>.wT=X���p�2��HxJ��������l d��܊h`�@A�nl�@|��[5��jػ�R�;Ul�7x�Z���ś�1{�^�z8FDNIg��DZ57�m}4��'�p���"��$�^���������O����(w!]��?.�00=�&�D�"Eϔ��fg��f]D��Cab?�B:�";�;bά�$���n�h?G�5��6Y/W ��K/1x-8�a�G��RbU|#>#��5���`��r�;%tICX��g�v���|��#U��[F����e�=ܿ}�a�e#Ȑȫ7FwE��u���#����I?���y%�H�Ќ�zDGǖ4<�fI/�/�.����쓰�az��=V�x&���m7Xb"���M���K�n�S
ad�o�L�����v�>2%�x&i�ͤb0�=���Y�������&��'t`����Մ����ʫ�Ei��h:I`7x�����e��z�����s̹"7z�Fϥ:4b��f������	�ṽo޶�/+�vۺ��\L%W�L�(6$x1��G��߇>&XM�Q	Xw� :*Zv=a�D���
��Ђ��0�4�h9������*G��{��[��$��dc��~��y�����:�O�aϜ���s�R��͘_��9��I��i
�f�O�y���A�y h��­��s����^P�@�\�m��\`gv7��ߡRxq8g{_�l�*���;�1�u,
�d�
�ֹk��@�kdj����Z�Q��
u�d �,���o����n���h���c��ʉ�9��]���͒<�ykK�U���!"a�/��F�7}����򣜉��7 &�&��򂝆;�Wg���l�J�ـ��IS<4���#W�Z����:�"d�P?�t\4���P;�ے��=�O�NAn�����e@�6����ol೬aD�N�oGo� Zc�c�TL���R��]�M8�-.ޯ���ű/���S$	�tAj[�!�����Dm�3:~�ep�kf�zmʀ�����|@�uX���	/��8�uŪ(����)8��W�I�/���Cr>��[mI�	�ʟ������"�Щg�pg��1�;��*��½/�;Le�6�w��!�8Yi��W���|0��d��;L��&�:y�5ʀ��d9W�׭�p���z�lg��q:�7؝�sq�7r{n���v�&)�'ޢV���K
��	'A�.hu�,��r�LjVs��or$s�']i��z��?5@�s2
�8���g�'*E�$8��!i/���D���%Y,-����#>�J�!V�<�<�~9����;%��P$��0��0��뭔�ݘ�R�K�L��cSx��+�5�}�(x��-��]�
1�4>������С�� ]�'?f����GQ��o�K���88����	q[Ѿ��+�����Q�.I�������mXo�h��T:�,�/ޒ�}T�S���
�!����V��~�[��f֧h�j%s���Ͱ��w1�8�|(���@pHlD%��c"�;F�W6��t@�Y��%�������+�1�~�^W�-����.0n���g��r`4�'G����俱��X(�/)B�K֔#���V&J0f4����6�m��r7Mn�&��������b��x�8��������ٻ�ژ��⸢������f�I&o�T�j���WamJZ�*�4͕
��-���p�Px�����!���(���$c��9���0 �B�Of;���	�s�W�^ &�l�s[2w�\Yq�b�%�|g�8���CU�alX�}I��;
�'�:h��ߦhW�Tb:n�GAh��/i��8��2#|D��9�m����|�A䕎�OS-*R����:PG��G�����yR���"1�=��8��͐l�r��dv�OZ�g�P��Ɲ<�h���U�o�7?ڹ�v���࣓Gi����xEHS<a���w�w�Ldz��9�/Y.��YHin]���28N괸d�yٌ��R[m·GG��c=�
����l���^7`�G=-��m�*>x��-��zv&�QC���N�:�#N'!����?��@eg����=����3G�L�k#�Ų-§��n�#&ۨ�]"W����VD�vʨE���Ӗ�ؓ6�����g��W��\���z:˒�\��u�d���om�_���* ����=fA�������� e�-HUs|H�,��@B1����@e}�?�Tԭ`&A�A�j�?֯�EB��2�w|f
�y��ɷQ��M���ǶG�U9�;�q
�d���a��F$����{����J�K�����(�wsQ��f�;��6UK����B�9u�T�)�KŽG�O�웃��{�h�ͣ�E��IJ�I���ӤY/�����D��#q��A�G� Y��v��DJ|��!�{q6�����o�h'�I]��`�|s��1�DU��"�N��j��P��]�,�P`�/k�\龇uJ�!�z��0,&��#�&rp[G��v0��>]�� (�==~y��C.�f��ؖ�I6z ���-xyb�ƎaT������IG�-�%��&&��)��HѪ�q���,'�Do�!���{o��R[Fk��6j�?�q���A�7~\�
�R5��v�4����IU��#5f~�~5c��s�0���� i$yjh�Y�&�9�Ǽ�F�^���b֢V]�L0릴p��Ϲ�i4�6��'�{�W���pM�9׽�ex4'c��I�T�\��FQ��K�t�h=@2�р�b`�����X�����?�<� =+��WH�ޟ�G��p�Y@�ǣ~ nҼ�q���ٌ�&���l�N�,�߲���I��.�gO���bw���Ÿ�3�L}��Ji,N�0��x���E��_#��=YW����t�-'/��|�d{�����f��������/�P�W)X�v:VT����
H4�5s,?�i��`�k�vJ���,G� A���a ���uSňB�������$?�D6�AC�Lb�Ca�s������%��F�Ȧ)J&B��ROK������+h`^���K�P'G-v��t]- C��=3D��&�q��/�m���A�@j�`��.2�Hh>��U7�0c��*���Z�l���'��_p���7:r@���䖪աA_���w�����_� i�_1P'/q�k�6����(��<-�J 9@�W&b��1e��;�X�nZ`��6�H3�&�D'�:�nX���b�z�Ri��Dܖ���961�+<B��n���H/ו�*����('�6��������캠U�١Zqqk�X}�C�i��X[O4��]�':g��`[�S�2'1�b
dC&�������1,��cW��OUv���7<X0��DPF-;�X�s��t!���S9��Mϲ����]v?vב�	?:��{�4,o�x����%#�e�08���G��q]���D���`� HQ4�"�ȁ
S�-K�em� P��|� }��q8�5
[��z�.��.�P�������8C�����ЎAB~��+�  �-��vE{�ԙD����d%�~`)��1�� f��L��.���I�/�,��黿f���{��g�^,�ͯ�T7�[�J_���S[�u�;�ᘹ�t��3�%fa�m\RN�6�9��ݞ�+�$�<-!$�CZ�� �U��g`�xO�!SE�H��gܙ���n��Z�Rl�ʨh��D	�P�&��Q٭a%`똝���_��U��\c��k�7��GU�z����p�� ��;}ύ��z�|mb������;H�H
x��U�T��Bz��/O���pzLM#"3}%T
d��Y�������T͈7�%e��B���uK��!�D�l�*�i��A7�&6ʵ#��	����<��XϘ|���8�"_N_K�&�*�u��v��oF�(Y�CO��`�jE� 4�/�U�ڑ���c�P�����8��E�j�+{�r���G�L�gZC�,!x�Q�P���+(A �Q#��\�r�V榔��?X*L�+�����أ�.6�C�/�Dy��<H���=pЍ��MP�0-yX�+�]��𲶁�4ˈ�&�)G���Ϫ�k;~�y������������[��n�����U�{yeQ��z���֜�T�	/�)$�77���v"��?o�$���3��G��6��|vD/]Z��K�I-z��K~@~�Yf�I1\Y�g��ه�th�C�^Rd��Ԏ�Q2���(�����򾈨���yU���7U�����Y����]��߭�pxE�'�6��x��`��`σwU�}���_�65�^<O$@�S������ƗO >���%/U�o�6~����d��G���4�(���~�fu��V%iu�K���8�O�0�Q�`I`�y~V���//w�-Ӯ�y2����n�\�P��7����+��썅�,���f2U(�i�v*� ˊΨ @�{^髲z*쉀|�}Қ�
����/K�y��y9��k]D�,�
�������S�����6m�t;��ԡEa
P�8��U��=99��9�����*�G0�$]1����m��h&�C�y�C�om�A�͌�Ae���_8��+�t�KYv<}��'�	�.Mj{d��"��@�0��9Ps���1�����D�	��nUr!��sV�Ɍ\� Q>�$ee�{w�B�D�t���0�:G��Y?��]�F�,N���d��=9�?7Vtb���)ۑ}��I�P�nI�r���)�uI �c���G�P�͵!I��\�@�κ�%c�1��t��x�g�X�+7���Wp���$K,q�Z����f��2�M>���U:�wR��w��:!I`F��$�N���z���\Ԗs��M�;�iT^U砤ȷV�:��v�SLSWb����$�>_��a���qf��5؃t�Ȃ+��)��~ֽ��Vv��8cG�U��W��8w��\�9�ͅ�n�����������#՚��3�6��9�CjHpKB@D�V�6�H���
e����op��BF&q�R�3>��x�
�h�#���zln2z���?A4�iO�#~�eM��n��Db��x���m��g8�3�(+şהiL�N´;ڞ�'�V��Iq\�����T��|�2O�v�&�_���W�iL��J�ޫ��JJ���Y�^o�y\�c����[�UH�(^4�l��m����{n�7�, &���a �sXKRtK7MHR�T8�;%����}l�/�y���In�0ė̬TȾ�`oZ6�L�OJ����膣��'���t����"�2����iB�)[���|��0:.�B-оU���D��xóo��ا���.���{�z����?���R����Z40p� ��w�O<!F,��}K��H9�� v"<����9RF��f������'�����{�<����[pK�$J�5�\�!�a��ݍ�ɒ�3�9���q�Z�?�ڻ�%��M�Nu��v����q�G'*�RA�MNE�(-��?Y�����Mo�:l��.�?���ݫ���5X/��+���b<�jV��z0?��%��uр
KH[�6�`춸�7���IZ<����`�w+b