��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����Y_��F��tw�p�^�=�����DW!of�.��"�"V�8��Ua}W#R�M�-Q�xq��ų�����#k_Q��?���B8I��c��l��{ͪNȽ�D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����~�Yp����ƄνC~�A��;�`�m�ѳu�0��9�c��F�B#%U����a�&���*.4��0�t�q��Y�؇i�o��!����A��rT�B.���,{��TX:.	��?���h��h���L�*�v�H�cO�(��<M߾!��q
vE�Ӹ�]5�����f�9� ���y��bи�{K|]6l�c���R;~����u}U���^��"zCqz.H7��W�u��K-{R��C�������D�aja���/�;�5�*��8�Ѯͮm��;$M�VEf�V��`C�y�l���W*XtN�AF+A�J�Jd;	�V6�mؤ�����W�!u!ߓ�~]�M����!h�����n'�8�	��U�YZu}��h(�E�+�lj�녾���&h����{��`|�`5#���sX��5�x�U
k���/|�*��ɱ,Zlߜ�S�M{�ģ�����X�KO5���X�;(2��
�ؘ���W�^G`8y���|�$�[��l����H�E�):X����uu�����@�?���T^!�}��c�/��AX�NU�r�N���BS�}��������Y����}{5�g�¾5���t��F_�>�?����V� 8�P��~����X�s�6��P��?���4v�_�-ֱ� ����Cܿh	��\* o5מ�Δw:�3�*���D�\1h��n<BE��z�ZV񤞁AL腋	O,'��R�G��ƨZ^:V O��Ӣl��#*&��/�����7^E�n�V{aߑ����8�go���@Wd�]�\�f�^��֢������${32R�|,"�t��u�)�;L`n�B8����tz{4S~Cf{�S"G5\w0[G!~~�J�{��Ұ�l�7��9/�6��߻M \5��5���|$Ֆ�N݉�8x��p�A]�/s9�2�pBetϦ=7��ɤSl�iB�+<��_�Ϻ�n3홭5E�ӞB��Ȋ��h{��h +���)�dp�Ȣ�1����ČET��N�d��nIo�LV¨Ri��a-V��5&Éq����8|��e����;�ͼ�
ZXa�1�d/�stmq�V���14���<�[�?�B
4���C]�N�(J�Lȍ_s��o�M�d�.z���#�1����{!�Ga��g�m�M�`��s,���>L�b���89�wX����,A dir_�L�&M���
�)�c�p�xz��`N�L;�7�B���_ag�e����L����1�i�|W�+��Q�v�D���MFߠ�L�9F��I�`*�T������Yʒz��$��]o��P�51��CQ����?��^�]����"Ľ��A�VQ�\��䗶˅Q�SF���q1��l;�u4�� �^nH�y�:f�1QҌ�΄n.*}Eu�����b���j�߀<��N����@KX@6A�q���;$9G]�4G��?2{�V�F(^��w��|����d���9������#�9r��/i�*FwC��<U�܊C	8[�T҂�l�Z�\���q�}�����u�����̈́��}�k��ʉ{��@�L6�YċkH�R�j��� :�&(����R�R�:�u�9�g�`�6�]���ȗ���+���{�ӵ�B�u�~®ƒ�G?���	�J������̚|٥'�A�J �R���)p��|�|�T���p�{��=
i��=#�?��6~��|�Q��n�OI"pE�^��{��)+XQ�N���0����ZNl�p�����w��4l�6=�a�1K�{T�@gv��c;��3��Z��]�����!լ������?|�xg�,�&��!<�(,�d6�떪H����`}�.M��CD�?Q�A�� U_
t�h�sU3%���_������pt�����q�o
��Q����1�-�s�B3a&�K�O�Ә��X
l�Q���ۇ?�!����f�$7�}��'L1��'B��~ƿk���F!��D���>k�2�g*���7\i��w�_K�	{��h�2p�Z/>�|�uG�B��1��Ȥ
�Rh%I������B0�ƕ�!N$\�w�Ո��R�<��I�;�����Na�V���ʡL�q��A��yN!�m7p�7�ZjFv	3������F�HW����1�Ԏ���4+?��d;f���X�t�{c�1���Y߁�݉Z
���:f�FO�
��\b=~�D�1y���ߡ�_ �.��Y��̏+j^go���|�S6(�iԉv� elu2��PK��=��P<�E.pqj�)'�Bf��ث+�8����%ψ��f&_b�ݩ���zdr�=�g�7}�񋏽"��,�*�V�HD���H��<�)>8��ct7��xB���_���#]�C���YJ���w���U��R�����b���ˋ|� ������v��!U0�V���Z@Ū!�L�(��Z|A��b����Q���=.m�6�ٷ�����#%�g�H-�|�h��(<��fH���/d,�@%k���@���+��^����+*�됵3cߦ[�6?B�?ZF�C�[,U5	JB4x[O^]�(ni�G4�="��k(4K |�v�Xl�t����\���.�9���ti�u�����u�U<�R1O�DP�P7uT�O���x�6���u�vhsـ4	�����;��ɓ˛m�X�D9��MR�Ǧ��&hհy\3q�f�|��{F�T�"�7������sɤc��v�t��َb���L&�O�}��3b3�:t��O�s�Ϫ���S�=� i
�U{ґ=���w�����J����z�����y=�����	��\��Ù��"\���V��\UƎ�~k��έ�$-�}$������6֟$V/�t��^-7��zWJ������q�32��D[_�3qI[�3܆pM�ƦWâ�H�_-񁪬�pT�v�L�e�2�������gLFR>~�^/ tg%��X�����d3�E�AE�^�d���!m�A�x�1�j���b�_��C�3������O)����һ�p.�co����r�Lݴ ��!�E�Gκ5�J��]�5$�{�(��Z���(���3�j7�%���x�CxXT喺�J���+
f�t�$�CV�hCR=�g-��-���Q8)���0N����N,U���<�ձ��r/���.@{��3�+v�?[6#�_��{2�y��f	C=Z�XR���������TK}vkH�֊��c�A�%Z���5�������hg��9Q���X/Gь��XjCɤ�#�Р��ź<�� Bf[in����s�b�4�T�K6���	.E��A�5XP4F������Y��X�o���J�����;=*�E��թV"��U&��si��;�=1U��]"*��D]Ν�� ����8�`A�6q�N��|n��K=<P����8p�>�A��Œ��2���«ņ�t���z�`�3��3���;�����K�5Ep,x5��*ZzE�gz���W��{A�PY�K��Ě�بn/7�hBc	���(69#��+F� �b ����T��A}�8��]EI�$��u6�x\̔��!X��lf��a!&QȌ_&�W��	:w�^�k[b	�) љ�̇��쬀S�FDt,��O��ۅ�����%�������e�ʯy�D����!�LE�s����9��/ "��͛
iQ伓�V�ϧKð+��ʗ���2�w�)��)s?�uV�rF�A�(��VgE�a^2�%��ш4b�Y��J��2dE����/�M�+����$��
�_)��B�\���$���D�K��-1]u�.�$9D���Q�RN!�KޗK���}��;^��X7�L�>���LOn2�c�G���,7�0R�|��Aw��p����xbF��H��P�<T�00d	]�b�~��i�D�jC����˧䷴Hw��75��s�5SgT\�W�9h��~|1��zO�G�\��/���td�ά� 2�A�VS����:���5i굹�� ^^����hAuBj��c�� �����*�+O�*ڮŕ|"��?�i�2a����"�bOC_��&��r��^\dt��.��I�_��>��r�%͏q_t%0�L����	T)�ڔ>��.$o�Y�f��}�W��Ml�
��'0Y��[bbEa� O����"��Nu����,X����젟g�&J�m<��j��1��\24:�k����"���QCR�w7s��e!	���/X�
���'I C��
��㠨?�/њ����A�4��Jm����Z�9A���`��Q���no��u%'OXD�U#�{KO�� ����!f��TiԤ*Ɉ�Ж4�B�A�*2dZ�����9֬����G#p�>�/n�;1@���I�>�Xpm�n����Ey^�VL Y�����X��+�C-��n�c"L�:��̧p����ns�r��Ǖ;ʨ��/����*nu}n����>����Y�,�d�a�-����87[���� Ul!(Xc�kQp��q�}�xU$ [m�e�s�)�՛��r}���� |C2�)[X"�ꕋ���ۉ~Ebѧ���$�)w��K�5�s+�_'�5ۻ�>���������D\S�t��+Q� ��vI�/s�B����?�R�/��L��e�ۧ��g��?Ҿg��[�x�n�_��>��i�	���Bm�h��U�.�l�Q/�'���Wo�����`m���RH�n(���w?A��A*�����^e�,c3CJ��9U�������|�ɭ���
1�8פG�c��'�ז�=ȷ�ƏT}� ,T��ćVP��)��6�)���ni��a�ٜ���ҡ�C;�����)�8/ݱ{*ǴX�O��1��P0t�g�h�-Ϥ�f�@u�@|gB��G�B��y:�#�$�Kq��AX� z��H:�Z2���Ŋ�{b"�q����kb� ش?��E��y�/��>T�~�rL��1���]$t#�[Tx8�4:��
xs!�l�s,�2��3U���������J/�Ҁ��
j7Sȵ�R��D�-?j< G��h�Z{�>�E\d�׉�4}7/X}��HFC[�����/,����A����n+e�t��=�3��%*U�V�63oIm����/�%wI��0"FN#���*�t��8I=I�߬��	Rй��0�Mt�NY�To�ZK��	��@�k�����`���7��Ok!�z�76�h�Aa^.7R]U�NAa��D��CBC�{�����@R�E�n�':�g����ŧY��h�-j�\�h�c��� V������?���o��*j�]�.=C�x����Sш���dD��o��7��K�؀������?�0�,p
�1~B�ˢ�)��tV�/��*:nR|m�D���Քb�X�aJ��bqv�^��U�3;�~gyɧ�ƂݯCd�L^���m�j]�f\��Y.�^���	�70���J���k�C��,�8�R!��}`��B��+��w�訪VNS���/"�Ѩ�ہ��2�qF���w:gK0:Q�nUP��(!���I3Jݝ܇�al�Yk` ��D��ک���\y��0��sr�[�R���I��̐��疬�� �k��6"�4cI'K�)R��� �; 9�t��oE�^f�*� �̅+�6gR[It�)��J�����0��>r059&��Tӑ�:��A���Qq�@�ǋ`o=���c&�+�Ɲz�j��j��٨��R.7(� Dq�����0�ؑ2JJ�=$(Y������ܰ!4�YV�<e��W��:���ez(�`z��-(y��N|TW"/݆r[u���WA�j��|X���=xh��v�h7m���vFg�����0C˝VQp���'�}J��]�����j�z<�
Agҭ��o�m�ij����P,-�Z��e��������Ҷ�d�� ��5�3�G���HG�J4%i��{�=&,��m���jVd4�{��n�ԧI�PF#��$dvσ�&�3�ЯZv��I�)4�[�Z����&� -s��m{����J�
t�I�o�u�q�cѳ_�4�g�rT�t�� ���"��U$o�����sp1�蚒Љ<��֏��P2��<s���CU8"D�3셜[����V������.��sQKd���N���� (]�s��j� u+�DMz��I�"���t�(~�3������|����};+��&�Z��e���"�]A;�g���҃R��}Ʌ���X�а/�Ye�
6�Q��O��B����29��K}�-��G��/ΰi�ۀ���~��å�U�P���*�SxD����H	]�!(��EC��(S��� ��w�;�'�t�|�%�����"5�����M��/U ˎ�zja�� :�HJ�)���G��ܔD_"�y�(F�������i��xq�P~B��T߆|���	 ��E��g�CM~w�x_2��b�l��f�ppi��.�A�e����{"�-��O�[M?���}�u��*�^��r@Z���Oat?餲����n�d�����,�8��֭� eR���]�HcA$+#Ld�`;�PԩmT�~�3P ���|�ο�k+}{�t7��޼?���5�+��rK87��:A�5�kd��C�\/�_`��d�B$	���}�Tiӂ��ϲ���(~U��2^�:�h3����Y6e�4��3�L�Qe�"�I	|��/\w�,)kTv/&p�T"�s%@��Hn��lO4#Cf"��P˃A�@��&i,���VE�B��*�@��~(4��M[ǵ�
n���KDL��^��!:� ��X8
$n�M'��A��(�%�.��)��餳�q��K������4����m�Q�/G�C��X",y0�YƼ�k�B��~����^����E��$�:J���z����1�����Tׇ���񱎊��y/wuL�5�-�� �;�Vty]ȡ��G-94#�n�q���֤��[�1��1c"��N">��tO���@N���}���WY�nML�#Q�6��{����8t��RP�q��Xh9ɬ�f���b-�����(lF}��nɽ[�=�)�4Hiݴ����4Y����]���.6z�ϙUE�:Q/|����߁����B�r��7W�l'훥�P��I*d�a՚{ua�M�XE��)��j��A�h�7���l�c�r@4i:�<
�SG�>����7�w�g���!\� i�oZ�#��/�aA6�K��^�ƊZe��i����� ���EA.�z:�f����+{��,������`c����08�w�7ǅ�)�j����8s Y�1"�G+�q�������#��pI�c���@ȁ��t��ރp�K:�U�*��^������7E���Z5�c����ς���$`�2���lm}ء):[��Dp��޸��g+S!���.(�����3���#�b����ΰ�2�
`��;�>�g,}\�~��*�D�B*���Sa��z8XU��4��-Х��Y\SA���O�	j�n�e����Q��u����am�qkk��I��1�%�	JdoMb��n�Z�ʓ����D�U�>p�ߵ:�D�t �);��O.f�i���7�>8�Q�;h�6�:��K�S��*�8�����j��e��4�6}�%ߞwE�Q@��,н���fn\��C��0iLr��5��Sc��4˿�f�Q@k˓nԒ�~x%��ٯ�H��P4(�����2k���Z�D��j�XM�X��,2H�o�l���hQ��-���>�\�v�2Nn����w�d�@F��%7rY�$Fų)��eԤ�+�a�@�2r�:��L-.������PKE����L��7|�T�`��Y��@�T�>�zo *0��1Y�ǴT�Ϭ6�g� �h����.VlҴ!ˆ����W�~��o�4���yt���~�G�6�b�Q��X�d�e�mw�|�y4�36��ɧN��2��B���|�kzs�&c :���L���W,���/�.8�mm��~�X��$.��1���8!�5�ǩq�1�1ڮ�m�##�&�\A�
v���2�{&�C�֢�1̻�Ȭ=�.�sJg��q�a�ۋ�@`ȬRM�E'�y���K$x�=�lij
;����s)�8��q-�R���É�G
���o��:���Vg���ӟ�A�Hm������(ԑYw���Fh�����p��Q�fĂ�>�]����,Z!���dW$��
� X{o\F\�5��FF���PƢ��#�I���U�u�-�ܠ��jD���O=��Ę&��\��,cl�D|_�͘<|�l�����
J�H9�w��f�x��[ �H���	1Ĩ?��$3�>��٧5����