��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��)XS}�d�v��rfO|49�9|J&MB�����P��R�3
ax4aF>2R;�{�j�V��p3y߮?��F��F���;�:ȴ���՚�W��W�@w�Z���'�%����F߷f\��Tg�b��`�lj(k��J�g��U���5*H�'�ݒ[��&���i����B0��98��Nq�MP�����Jh��X���80���%�r��t 51�������I�ݢ2�DPCJθR�X1�ĵ{-��
�Sxb�G�ՕY.�CvG f5p5�{S&d�/��a|���ԧ��R�ZD����gu'>��U'��f����c�'���}�!���7�=M'"��W]1��Ƃ�͡2:��q[�R�C�5�:�T]�L2Ey���Ñ�[ғ�&�[�j=j/$%u*O |����t�&� T�in1O,f��@�#�����}y�_�[�6����EL����D��7�P��ݖyt\&T����jA���G����O��Tix����w���]#�7u�^��m<$֔<�Z-0ž�]EM�pY��oS����ǫc�n4���<;GX���樹�$����|���Q�s]��g���4<��,^� ��?�e�Ĭ�ʻ ����i���^	����K�#X��e���Pd�6�Z��Bj�������δ��\��#�˴/r�˨HK��S�!�A�*�L�8c��	��U�7E�Q�K������r�k�R�"��S���m�S$�^�I�����*��@w��ŋ"=%�u�� �\��k�DL��+5I�@uB��0If�#IGh|�dPV"�8�JT���y�_���\�[�D���̴�|