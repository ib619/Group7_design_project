��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`����|G��x>!�Ш~.X�6'��ӎb��:c��SqՉ\�Ѕݪ���@:�9��y.P!�O�R��F��e�:�G	R��H#� ;�ю�gT	���ݚԟ,�pGpި�W���$*|�߀��0V� �9�ھ�w������y���zNq=?���`аG�#(��.C�S���2��bƬ�>b�N�]{��ƻdˀ5R
Y!�������5�/rsK@�>��kp��]�K��>��k�{9�l;0���J��[�x|+&Lqew�:z8�����.����9�\��q�c@�C�_K$>Y����98eb$H�KSH"��Q�� |Қ�,�-��{h0C.��]? ����Ԅ�/e�w��i�����/g�CVAi�ܲ�u�c�\}�[��!��e�:vM��c���Dl|���f�!�^G@�V��:t��"%P��$+\�5A�8�rG�/���/�m��S�"��_����������DI$*T���F$�҇�� E���\�H�A�X&tI�W��4p\SM�S{�!
������ %��O��۸z�H*��1�A(w�A��d~(�����cf�Sp"�	�,4_׼x��\��݂�$`,�P]I���Ed�v�n�=���g�4o܄�j�UF$��y&����``�KRƓ��f���P�9P^��์v�L��Q	X�w��wYw:x�����{W������٩1Z�F �ě��������P��"�n��nj�z	zy�s������ІG���r���p�^-Pı���2�)�©k��n֥<�Y��f���J���'C��Q��.>��.
��V���V��V�����F�7ʂh#U��d����_�ZB)��JX��L�>S2���T�iǬ��]�<V.��	�U҅��&��fHz�![��5��'��YL-���m�Kɟ�ㄜ�L�߷jUΘ�Q|x��p�쬐Z�m\�f<�kZg��2"�F&9���	TM��ab37JB�b̔�_āWX$�-��P.Xȝ) �vO�̖UbUr�x�:铯�=����X1���=q�3�3L�E,��z��m�K��(L��
|
1U��Gz��:�ݤ��7�g2�����K��&NfLt�*��n^?�>��6z68���|��^JT��w��9�	2�"@���q?����c��q�9�a�nO���nv-a΃���{,�1I:8c�rf�|�mD��t�m����7feӪI[���?Ԅw9z���t�{�� �4=�2/΃�%�����E!�Ly���t��X~�&����<y�]��ŢJ��\�FuFܟ�ʠ�[��bt�E��c�h�C��@�z���So�	8�.T����j!��T6�k+�M��[9�lF3����Hҩe���>Jl�í�H�}f\���R��6�3W�j�j�J!EC�����Db�J�bg��7������d���8��Wdǀ˒' !�Ny�Y.bF3��R���dM`+� � ��:M��Bz%pj�.�oƉ����ߎ��6��}��Ӝ�>��*G��}�g�\ 6�*�y�o�������?#�<����h��&v����a�~�[@m�y�����Ǹ�7��.@�>�n�	)dT�U��L�?�3� ���N4�?����0œtX�2�J���)�k������n�a0a,��L# �b���w�̧^���ސRjY�!-3��G��g>X���2?#�~�Z������R1�\3H�&6�H����1�!��Z���Ù��r�i9�H9]\l�F���>LD׀��9d��{��+��:�6���D ��bC�w��6����.��p���>߂���*���A�����x����Ga����&��t P�îk,�vd��Jj���rZ#��q�����_����D��A�r�̵,>a��)Y��_�.��'��I�C�\alDE	vl��I�zI_C�?x~�$]�����(P]�k8K�d��Ow�?UQ�./���EہC*J��R.��UZ �]�w�U5�M���x��ԯL���q�4��x+2���6��>�G Я�e���H���m��)d/=��m��t���XiLfo��=E�*�z��"p��-q����$��:�����]���|71�>y�F�*5H�0$�2�������-��$���n��nU�f�,����5/?v�H�YKe���5�5RT�P��$�VЁ}���<�f�����4)�>-�5�*�Oާ�wJ���ALz��2E�x�[�yҊ��r�Y
�=�(�,$@�+B��M�|�/�T�zƞ��&�W�K��0c���\z�` 3+]Y�;h�s����+Qu�9I��H�Y0Rפ����ٙ9�w79}�ӏ�0���l-����t�R�z-vA�䳫�]�Uz=���ԿO�����sU!b��7Ǩ�I��2ڤZWK9~u�Z�T�l�n�2
$5��<-�$��R��L?��ߐ\G�λ��q�3Z΍�}���9�l?��Ü_�f'�x#'R�!'�{�~�$�Wˌ���ļ��3�H�aؑSA-���v�w�X��"x6Bc-���t�i�i��C畆���>\E�����@�g�v�	���{q `�xԱ��a8FK��Ҫ�U�Q7��.����O7�W�"�>�K*⌸gNR���>����k������+'Ѭ-�o����?~��h�E^X�ת���U;A|���)H�eflb("�W�]��7�Ck�.�������o;�O�Z�0�ΫkN&�<J�L�`�������)0
���WX��;�Ǵ�n7�F��(_U�u.ԍ�9�W �߄Gp��~�B����_P@Hӧ��N���AB:�|z��aA%�Q?5����v�a9��q���B�і�G)���6�6�ˑ0�<<cuw����F�9�E�V��L�)�V@b�3�my���+)�!p:������cC^���Úr��Sޥ��-�ӎ��;�l;f�/�G|.��baj�[V��p,�j���z$�V+��Bk=����6]-�$�v>���Qe�q�q뇝w4�C����ecO<d�Μ�\[���}���2c�pʓ�Y�lBvޣ�V��/?�:=O#o���)n�DI�0�`Lvt�W�ۺR�dǖReD�ќ��XM	^)�
=�o�l��@:�od��U�A%�lG�;�U� m�hk3�#[S�Z��<��E+P�.�BD	��oUa�����E�{����O�cxf���@j�ŭg��Cj9w��q0E�@q�p��>��X��"�6ls��AB��|��M�,�t���~/~�	In��I��7��� ��Ͳf��3�,o�0���0p�	�/|���`�P�ʃ�?�7���~C+v������6T>���lyі�ݐ@��r�r��[S�ÈZ����P�����G�/���K� LMy�g�,-��Y��𽙆�L�e�[O>4|MHZ�F*��II�
�n>�=Ӎ��m��Q���Y�np���hoÄcC��

^��t��m�3���IT�џ����T����ݮ���~� 7b���G�¼-B)A{v�@I0�8g��UI�6l@���C���=8Մ}���a���~r>�:�h�UƓ��w�e�(�ƽ������A��*�"�\�b5b�6=wd�T�V��*�a���Z-������<�)�bk�����o��v%���E~Sn��t
����zׯ7��}B:�D��(7��y�$��e锲����J)n�d��P������bօ?CB����ψ�p ��N)�8<4�J[ �Zb��c�Tk��dcr�7ݽ���^��g�^��g�o�Z��;5����Y�|�+T/c�0M��x��korm�j�V?�h�+�!��P�d���V�m7��[hO��&�6<۪�HK3��:�\�ǋHf>�s��Cf/�,��J����_�\�)�� 7��E��}v�Fwfu�x��i�:�n�BUi��@�p�iI��.��7�^js�F�vR�Y��q��sӲ��L��֗���bj:XJY���UD�][�o-ЌӒ����0.�Â��-;[��Gr�rU<�{�l�R�mLmo�,���;�z��޹G����X�f�tY@�3$��B���F��묛8�1�*>��B-C�v�����1<v�B� *�j/�?���̩�6|R\z���(<�'�M��^��/i�a�8�	m<=��X�yT��������^���\fiA�8TN��"�c�wW]�o4��o�zcߤ�� n��TԂL�r�N��6��<I?�_~ �U\:մNy$3􈺚�[]�
��$� �K(R����	|j�S�����iI�6�2qP�;z��X1SqT�_A8����e�y���yO�[5u���\2bXL#�H
 e�C��\ځ�)��jvj� �¨��7b���G�C�f�{N�EIeY��o���6I��V-xj�JI0��ɠ��˒ᬛ�S܃����?0m�jn\�l5_���F��	x���%V�C�k��`���r2��īV"R��k�|�ȵFh�ƥt������X�7�u�!̎�/�}�%
�����*�8���O�Pچo.��Y2Ԑ"z�\2`��?1'�5�Hz�V������Z���K�0x�}�w�,g���Q O�4o�:1ش"��xk!�N+�v̝��9eP=��>��3�V��d/����������W׹I�"�gB/)����h��@\aw�nFА��(VQ��fh}|���>�B��;q����fQ�V��qH&?@��K�*�\�K`c1�G&��Z��P������� w��1��Q-K���'�;��R��<%<o)\ �($G,b�b\6?H�fu?��~I��`�� $���x���
5�{���n�;�{� �*y�g��ۑҧ`��@n͊��C66��(Jr9T�x!8N$3��@W�9�12��ڄ	v����"�) K�s�M�@8P�DѰq���3��f�F�̞'�/eR��)�_L�loy�VR��{���24��{��	���FI%
H��$I&�$y���5%��ܪb_�<���ϖ�h�٩�lI�<}�'�-q�x����뽼G"Xt��ϙ�������D�D��\��֘T����"j7�Cݰи$�C�VmX�%8:�|}_c�39-���'y�yV̀�@ :��W����!��e'�{�s��Ib!{7}�a���4
p�����o�.g�"@��d�ҷE�]A��O�F��7�3�B��x%��-���#��>��:+�{H���o����hx����G���@eZ�xD�ӏS�������X7�7����|6	�� 2uq�Xl0����M��