��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����Y_��F��tw�p�^�=�����DW!of�.��"�"V�8��Ua}W#R�M�-Q�xq��ų�����#k_Q��?���B8I��c��l��{ͪNȽ�D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����~�Yp�����i�`��� �9�Ĭ�N�hh_��E�L�(�-z����/�I��l �J������TH��61Bl�J)��ɓ���_�Zn�-㙅N� ���je��)��)a]XOX�[:�"Ϝ�eq��S,2�@	��ݟ)\���{�
'�\O��j=w��t�e�D(�*��P����S��~�-2"�'�����FԢ�6]�V���aX[Z�(Z�w�ES�n�vq�#w�xEY��ڌ�(����_���PG���e���λ�9���9��s��է�j�Q���〝����uy�_���8�|�z����mP��ce����\��������	"Doj|X[a�)�. ϥ�ɉs��5�o��S�$1Őo�)�������y���⏟���r�sD�!�^��r���S�t�2|���e����������n 5T�ܥ�Qѵ�IeE�����}��+�n�e����K`�K��w�c��r����挳�s^�Vu�$��@6/Ne�m�AchS��}
�__�׼��4=����4Υ�Z�\T�� ���$W��M�^���+�0��v�~��;9�TD(�AyL�0�qn'��P��-��^7e�2�m�^�,dp���%p�RF�R���Ay�h��P��e���#'J�Ș^}�=�b�Z~���NԕP�~J�).n��+�t*x%�N��������۪�2�����ԝ�E���O���,����L�wt@���@�����$��Ң,A;�9�μ��)4a��v��vǩ�{��3w�)t�WX�R5:�x�z�)!�'�c/Yَ���[=�毙��W���h�PŨ�+4����2�r�S7�=~�惞 ���[X��*d�u���_��$r�Ѣ0�_9
M�g!9IE�h��z�����)5 �'�+��[��g���6�7�l�M�/ߪ�p�u�k��
��7%r�OF��k�[�r�͉��s!o��#�q���̖P�������5��l�=�W�3�p��lƷI}_{[e����� 듪s���,Va�	���D���I<���PM�w��b�T���������ɏ?�hh��Δ����E��5q���q��&����@ev�U��ʕ�áa��e�����/K��,�9X�=u���C����<��
k�d8�雿�>�1�1~c��	�jh���uF5��ꮟ���{ls����Wi�r�j��x��_JC��1�9x�06rN��]�$��_�?�U�˔ɇ���;S�zB%'�Z�O��a��N�q���� ���%_�|a��hCV��r;s(��cwᷯ�F����2�7�^< �&�7�j3��zf����u/�::``�x���$�dN�Z{��*�OwG���o&��LS�jf�jH
"���o���+��w+�0�h#���]�x��ʺg�h�7�`wZ�H�D0��N�2���Jf�H{��:��I��A�;�>�'+=V��]FN�06-��/{�B?y�J}c0�S�����C@Z��g�����J艆��D��À���x|i@�Q1�:����$HF�\L��_,"8ݬA��nه�����5x�XL�M�As.��|��d��T�a��n3|ňܪ��C<Q��t)��e��$�DzI��2܎�$�����P�W����e�=�U`ѱE��m��<��"
��ȷ�G��6�}Oy�}�Q���ILpa��L�e2Pp��!jU�βr��%��u�Q��7*�> �׏*A�(���y�x�ǎ�r�ퟥ���W�ݛo��/�����H�eF'�w.g�Qg��S�bT�?�RX��_6y���	�q��5F�_��d�x�3.}|O��K}�d��W	��I<t���A��+ʩM�\�$}\1B�(�
n=b �%c��=9Jcb�/n�������"��y@oe�/n��A�7ݨl���ؤ�e=?���'��#�@����9=z3�_^ �yDe��O��%�j;RmD���O�KΨm�g�Wyw�A1�)���j)"��]�g�p4/\"v�sg��~
�������g�&�ڥ�ʭG�[�Rg�G"Q����SK]9��~
��y3
�?
j��.O�v �v�>F�k�gl�6��'jF��=�Zid�_����g���O��i�fKnϧWA"�5>��xT'r��=%�<mK���OϮJ�ں%���P���F�f��G4��y�'���\r0}�����!Y����[�O{_���߈�Z��#�o����ki�����V���nd��<+S���Tt�BhQ�<8$��EҤaBa��]@Sρ%@n��
�{OӃ�Z0��lUK�C8D����c )u�T��d�:�J��)�^�z�%'����e��4��UI��W��:�T\�ȧK�ާ*>����ֱ����z�b���a��*3]:�s��HT��Z_�T��[���.#cP�-�V��-H��#A�������o���'k	馝�
�/j�S>ۀ�8<ܣ��"I]}!����=�M�3���[O��-��zB�<�)"��MQ�Z�W�RuҾ�ގ�)��v�tk���lt�g�Ki�������Tv��/�<�n����'a���)=����k}Ɇ��y{�sa}J�L�Z>�&a|VZ�nR�^߆ot�1�tA��A$�0p<LD�*���&S?�s��Z2��x��-`�p��f�s`�3%�:��\e�O��B�r1Ja���g˴�DC�+�p׳�>�ÊU��E|@�kX@0�Ѱ���<���M���v� �٘��7�;��m(�w��Es��v�g��&���+?J+��⌗ ���`�	 W21���7�N[���K�4�ۛ�����h|�M�������������|�V�1&ĕ��X���4 ��$�7@Cqs����K�ns��9o;��;umL�_�k���^w����P�FÌ����|AW��d+��B�˅��r ��M����%��ޢ�����2�5*��������;,m'��&�v�Жt`�w;�#pC�$��tj\i׳����D*ըo1�2�<����~#��!�~����,kRb��_���sq�'"nviGy��O���Z##�=�r�t��������=�6垵�������I������|���&=��|L�iQ�de�z�F#\?�|�@M����eN���o�t�We5hL.L%�\�ټ�l#�YS�l�F�]j*��=����z|U���a�6���g<�]	�"On�J�(� #����t,�^w�A�ĐC�Oㅎj�J:� /	��	��{�?絹��u�ŕW#_�{ED�/���!&����!�ֵq�d_�h�e ���-]���ɶ1[��-�ꩩH�7�ns���T���U�s ҽ�~�s��Нq;�@��-�|������|Fjϒ����2oP*OPv�����������C�T������N��.;,���b7�ç��L� ��GN��Ls��9�I��`�Hxg�\�쓐��W4�~UZ�:�#t�՚F=��F���>�D��Xp�4�n�B5v�����l���<��٢	�ds�	��8)b���u����ϰ�!���*��O�mj�X
'R�w��	��_��sM�#�tP�ĥ���w�ϏQ��}�,1��c����f�!�Cdq�je��Xn����ʲ�0���q�ּ~᣷���$�Yp�z
onQ	��^�&�E`^ߤ;��,I� nb�9�I6�>����Z	���ҁ45�����0w�F!!��+����~�ns�l1��KG,��g�+�H�v��ie��0���z�RnAw���4���e������qد��,��cn�B�����
�#ڈ^M\V�\u:%�gq�p鳬t�����#6��=h��VfW2F�Blnˣ�e�����t�MPm��<�� ��'U���WS&|��|����FAv7���h��<G�x2XC��ds�C�ׯ1�V0.%ӟ�Shrt�H~��'нU��R�
��4$�Ɓ*%���U?b�U�}�Wq,�/�.码����%�V$X�A���K�VY��z3�R�*��1�؂���7F�b  oM+�M�[f���P�	Pk`^����ۃE�5$!�F�)�B��L�&�d<C&5]`�% )$�,Y�W���w����IF�y�]�7<�xķ2�Gd:��TG������L")B�Z?j��ڊ�]'�=e�Ԫ,�/��@���|U����Y����X���a٥<Ri1��P�����{�ϓ:��`z�LZ)����|�b��ü�����[62���PH���ΔW�FM�����0<�Z�7z͠�8��<Y�-5f��f<x��Ƥ���ɟ�[J1��cVAi/�c�!3�X\ 1������b�^U �+��׉�q��Z��%��q�"��PsB��t]��]
hc?�ӭF�FL��Ҍ ��t�A�ɵ<�����w2z��E3.mq����	��s��q�і��7��}<m�r+1��at�Ӱd�`eǭ2�S��X��p<T�;�$��J�S�j�O���"U�2�;�������,(�=�l�����w��j=��9�.�He�қ	M��{�~��?w�f�'l �?����Rz���A���!��O���ք�^�񬞪tn5j�"�j�"�}�"����?�IR
�;J���Z�q2��QN�'С�A�8�����"-���J ����e�n`XI�B/b��\�pUֱ�ŝs����;��Y+Y�t��T��xm����9�"<#L3%N����J9� {/@me��&�ވK����w-Rq�$Sr|�ӿ��!)h��� T�z1�����k|��������q^�/�H%Q��s0t}��[�W��B!�Nx���Z�
�׍-1@U����ݭ#��tn52`P&�!��
41ޟ��A�`Y	�� 4�sw��zh�R׮��	�]�5�f�޷�)�©N%X����=�BGfB�	p���@��:1��.�@�O����(:��{�ˋh��f�h)*x��ݶ}�^��	y1�8�:�5��zAx�Řh4U�{z��`=���H���7���_n^1���q���
/�5��;���<��<�(I���&�G����|s�ID�H����T�L/(�%[���e�˖R�ۆ�m#�)#�z`�x}}d+"jѢ���`��x^���#�0���]#����7b�eY���/��w��F� 	�h�Ї��_+M_i���-'M�@Э�Gߙ?C���tr�J�y��c,�ǥJOUp�)�թ�r���.���R<�J���y���oC��Բ�y�E�}�,��).HR �h������/��-E���V���
�x?�XTS.6`2(��~P���'6(��K����~�;�a�1�<�6W��,ݖ�cnu^�dJ�>��\`v^�D�DI�.�FK�������ެ�?�F��VL{<z��׵�3M�W��M����<Z��7�r���Q�:z^#��ٚ��aO^KL��.��0.Au���6���U��J~u�m���|Ԃ�G���pܴ�X ��7�<����=�,T7ib���8j�n�4��J(��z�]V��^86X�W�������s�V��^?��K���	�.f�+Ӳ��6�9������b�'g�<č�hR���&JK�E��u����shB�Ʃ�g����Q�[��n��W|���C�~�'|Q3u��y��t�{?`D�_�quYw7"��1!����e�k������foH���#���Qw[1�G����j.�0� ��<�w�K�,>����%�F�W`�{ODJ�iה�N������G����C�a	�ݺ}�X7���d?r�@u'�<YH{���/Ol�U} �H�[�
�j	���N�?����&,��7)�}��uSy����e�~����݀_^�غ���DgD4�4�,Q`����.�}փ�t�R_����*o�6��hһ�"�G���Q޵C�"^:Q4��a�[����ᘍ�΄#�1�������k�c�"#�������d�~G=3��4�~wy=,�l�S�ᛯC�U&A��=C��A��P���g�H��W�'�Ƅ\�ڑ t&�r���m�����2���6�5���T���K�3��bg��D�u��}��T�6&V
��rIZ,�s6�d͎�mZJ���Q�D����C��mx��3|.�= 6��Ax9ƂM��+:MO��!)	��hrn���e/Rȳ��ծ�v�_]��xj��^	ދf8$9���ؕ<��MAab�e:��d-�Z�{̄���\��ߚk�f�v�ژY�k���>@XF7�3])�gD��'�5��Y�c����q"���;��`��N��C�݀�e1x��P`�X��Ώ�=�8W0�`<��S)�.�h���5�W���>�z����.��4Ilp��s	����]��Ώ,�
�B��ɂl�Xr�	��~^_��Y�{��0���s9eO��^8�>�
����8�X�nܳ����@�o��	�S~b�Vn I՗�O����M~\�.��A�e/��vN̷���V�?4.��J�2\���u,��kd�=���qq���2q׻$�_>z9�jт�� O��蠘Vk���f
/
y3>����Q�����r��Z�
?h�K��"g:8��,�-?��8�T�3ըNj3 
a��RX�-s���|�E���K��n�OQ�R/_A��� �p2�S�,�t.��Ox�7-��\1�����E�iʨ�S"P<O�i���}cOR�6R��bSYW}���뗝t����7��#�g�ִ]�J��b�f�ﶝ���9��1M����T���PѤ�����;�R����&��<�����(�G��A���l�w�M��Z)���uS䔢J��\O��ȅ��0�����l2D~􊩻�`�1�r
��NNL�ZB{=� $g�9�d0?]7 �M��}S�`��Ô2���mr.K&� /����7�7�ҁ{��ۓ��9d���e.�'�(��ŪcQ^���g�l�G4Ѷ���÷�j�Q#"Oȱ��e,�yI���'����_\�|�1�A��t;b��Ɗ�����)�4�Q�ȁ"'���[8��HE%8���/���G|)������s���nĂh�.鳂Zr(��U�JNv�_�o���2z�\kiM�{��Rq~Spl�9���Y���"r/�������Pe�!��&��B��v����w�`{����  }o�X��zC�_"�O�H��Ҁ@Ĳ���+i=���������O��k����OT$r CVy�m��eA(�Q����-K��iv����
t�ŷp���~���z7ޜ��5�>��KH�]�����L
2):����h%0H�3^`~�{Q�z��9�|X�J1M�
up�~e��+�Ц����5�^�)�N�탐���[��Q�%qz��w�v��&�p�^
 p:�i�->eg-K .��c�n~��=7�cՈ!��V
�$�~�2�ZMߓ��Ԛ������0X���q ���3-<<V9�<wl)ag=�s}F S~l��ز��h�_����g��~twms�i �&i���1��o����4�*i�2�D��%f�D]*�^�P!g�(=���
1��/���|�c%�]�S�l?��G����m��Q��	&�=�S�����3���cz��Eh��O<kcwe����哴0CL�⨫k�u�6�����=ᗐ�ƨ=H��buM�+���J��?J(��']P�V���}�L�C��~dM #�Yۂ����?���,��'j��&#��O�-0U��l*��a��2�nݕ�wiFl���E���ɮ-�k[n]������ v�;��Ԣ����>���?ាh}%����SS�+����)B=�O����m�G��9˺��ڦ4J@�(�2��y�&�A��A���Z�%�n)�YY���`f���C�;i��C�=��i2�i\��b��f7-�����+�e��=lv� H��DX=��{�PA,�C]�d���;�+�5g�T��������V�k���/Vv�^@t3u�F�E<]F��[�*b�zR��7Ms����32��i�sh�ECll�hZ`+Z)ᬐ��v&cAi� �3P'�5D=[R� ���+��*z����H`}$ �*W�#og���d69q�3v�n+<O��/B�-(R�@�J�9����l�k����&B�k)w�B�<UZx�xIS�O�v#+/I�Q��l�4W��Az�w_��I�	oP{�
�Jѳ8�_���68�[������:��Y,t��׌��X�Wvx9��$�~�Y`�	l�v��l'��>YI�dY1���?C��.1f�ed�R8f�xwdz��S�U�oj�ҭ\��/
w��5�C"&Q�ז>G����Xe&M�����C7rʍۻ��SI:��FbE�z����[�'3�}��D�빫�5v��]�����M�k�vU2�<j�jK�2�n��b�i`ɪ�8�R�`�ǋ$�j{)��hl~�bȼ3Be��t�����,��I��{L2�,[�}_$�|�&���L���v��l筻��..��uam�#��M�x�[{��P%�!��d�
��@F��=�ȍ��Ik�
�]����~�Bu�� ���؂�G�l�C��7��u�tU=�J�V\T�B����~�����9蕛 B���][���ȷ�F͊,�;�W�3���9iܠ��?	&r�K��H�`j�d̐E�CP+��u�����0��c�UU/��Ż�׶�k��.+����,�D} �|8�,"��j�]��h���Q`��i�����ىzC�Sб����Ϫ���s��������\����� ��}u16k8������l�7ܓ=_��4�� ��&IJ�a��ΰ��`�6/�$+�Ńɝ��L��J���	0�b�Ei�h?�(�GG�L�M��Y`�I���L���O��.�f��
�B�f��OȘ�h3ƙɾ�+ƣ�X�%	��p`�p���@2!<)E#5��8�K�؊�u�S�i��e*3!�d��N�	�$I$���잟�ԕP�{~�Mu��0��WF|�& ���o��N�3�ϭo�chm�5����*���K&�߂Y׷%D��N�%\U&*�Cdpɧ��s�{3��n�VmP�C�I@w{��Lb։	iW�/fU5
	��S��H�O\�Q���zsdJ �y�#�f��m��Ks1o��k��#J �V�W9�|����0u�'o��ݫ�F��I:�EX/I�Z��mN�<3i��P*	�-�t��.�`{��m{O�l�ΥHko�<�����:�
�b|S�9ܻ~3�x�s��9e���:$��7�ZH�2s'����4�[�"��i6(?�ǜ��c��Si�t��	sz��H�5=]���Y^��}���:�G��K���t���P]�������FG
H��	/���ӊ7]/ep�xh���h�W9g��g�cT� ^|u2缨�;��+Z�R؎�:^񳊗�Һ}�w��F�;e`�E�m��'���E�:�f��fm�0�R����۲K�Gm��^t����x�=����e�`{wEDH1.�z�@�~����E�;IO R�d�Mu��<��#�K)�;��	�3�+�<�P�;��zwN��_5��4�=�U��C���қ<�����iT�����?���><�Ci�R�������į�-	�'cJ�������b��M���=��c�+xI�Q07���82N��>��tK
潘x��w��۫�X\��	.6\�rC�sg��'�)�-�,@����3���2��7�j��HГ�摕��;��b�j圉�7.f��Q�Ç��o��z[��z,{�R����7��#	��@�,B��E�(s���7?���*�K��H �`��wљ��E<��$>��ʦ�dAX�"8�R��'��?��$���"f*D��E�Ob�:( J��^��ʧL�U��dw�I,�-{LO�
V�6���.�>��[㼟��p�&:�	�t�՗���-�ť^���&N"Ʀ�jD��ݠ��j�m�X�]�n�
x�B���W��19k{� ����G��ꈂ���\��`I"��-`�f�Z��1��=��Z�5�Q�.y�yN}:��| Ho���/]�ԇ�/�af:Q�O��1D
6O�#��n�A$*���a�w�.��ڹ�xP����R��A���5��E([P#'��TRG�b�}� �UQ����|�W�����y����t� �V>+���%Ҥ����������`g�^\��^��.�:��Ha�)%*�s�[�wCi�t��
[��pe��Yw��PK�N�f�JS�ݞB��# �V�$�V.�KI3|R]Њ�a!a�ς	Ax\����Q���y�#�"��FR���!��^���]k�Ňmeɥh(w�Id��������E� 47&�T�2���!���F�l��Ϋ����v43e�ݕf7���BwJm`&�o�1�� I�=�S�����qh2勓��xH����_!��w�����F����A0{�p9X«�Tց��JYw�����Ĺ�7}.B�Ú������ڝ����m��>�^їP��3a��mjč ��|�	�>�^l4^|%	���Xޓ=�lSO�8����-��HR��~�TFo?~�HL�!aXW��"a�6&_��9.�:LV=.�?��%�3�aQ��wQ��B1�k��=6�ػX�b�uD'���*�H�����5�I�3��Z�`��\���6Q���QY��
����;;��:{�2���C��(�wM��ޘ�w��KT\"��J�F�&�PX��)�Z1�a�7@2n�� 
�$����5Y{u0Wp��egW�3�H,kr�t
��wU���_�Qʍ��_��v??gĊ6��R�N[�|un6V\��ᄇ������`LꏁP����Q1�C����$Q[eoi�p�co�BQ1_/��MS/ku�~��P2u�8�u���J�&3�0� �
�|�<�e�&H>9��o$�\c�e@�����ڣH=\�#/Wd�]�;a��������<
c�|!�R[4��q.5|Pm�Ú4��L�V_��`9�*�@ ps骥&w:��,t�>KJ�i)G�1ݰ�J�v�"��BR�
 hPA�׃��������/�\�n���C6vl\��#�*��8�3�=���1��A	E-�E�ܨ��Jl���l��6�xe��;��\�������������  E��\���@����!ф๘!c�ƶ���a] B��O�Bx(2�<���5Kֈ�E����2�m�wJ}o8H�:`��H�,���˻dy�W���� d����ʋ�B�+M�Cv�.?
��6\�^ٷ�٦����=��L�AK$��q���sg�����J���@h�1��>���ogǮ��?,�(���!^�-A=��o�Q?c��w~g�-�T�nL�>�c�����!��,� �	��1�d�\䳋�=Z��O
�(ȿA��.ʖ��:|Qߝ��7c���(�i�47N0j01�i��|�H0�̸SR�� �/��v)-�V�%�#����W���rПԤ����bˍ�)�#@�L֯�D�&����n0�5��[E&m�7z���g���@�Z�j>Iq��6��t��ŭ��z�.���3}�Fo��)�>�ϵ���*G�����|�EykS�Z����%�;?�B�AxR��ay�XEerS3�p�{�e2�f9Q;�z%N�v~�g�F�{|�l����K�Q�W�߹,sҬJ�Tlw[�{�kx��0h<{Ve���[0�Lȋ�3�R�A+�������q$������a.3c6b~��mk�?֒�>l},dD7��)����M�D��j�R�2��(eB/�tL� ���8�{:La��֛"����=�l���{��=�ųD��Y��W�p�.C��nf��E�l��(�5�o$u���A!�+�~C���Λ��3�%T1��fH�c�m6p�:�vPi���v��Z[��{P��7�x�ix~T�rN�)���7hf�pKr�6�=,.<F�!��*�P߅x��Le���<�5�gk���Srr���Nm�f��Ń��cl��Ή�V�*�=_�^l��êa�q�'�@؄��(�YL)2���kF9�ͮ�����q�+H>�H�v(o�P���b?���h��l�v%����n�����e�GyB��[Y+�R��Ak�U���f=���&���^T�L0/�6��⮤̂�}P��,q�6�*KAǧ'I�!���"2�4�7� J��P-��FG��'j㸌�m  ��Řuj�>�9��H0��}���~��=�U�`�.�/p�-���R�cm}Q�.��6�J�����)vSwѻ�XK۶~�I[l<nݴ8f(ɰec(�����dl���/��+��A?>�/H�
�N�-�6�N=*ml*��u�-\I��D*}{;e���o���d��Wǁ'�!8�̺�l���MB{� a4�c��DImpC�e�ӹF�v����=!��8 N5B�ک����%���ۭ��e�?a��|Kq���Y�@_��oܵ�r����A�'�V��/j��l��aa�����ˬ��GM2����]�&�^n!���:,ȐE�b֌L���<��Q���1����]/
{��V���ݴKe͇��!�����kn�W�Yq����ա�)���zV58`��:���f��2v@[b�u��H�3l=ӿ}|4�C`�"T��gE5)G���a��������T�~�D��=ɞ���B�n��R�oΣ���wK��m.K����J�`KT�����H�Ψ.4>�>4]�����s�38�aP��0=*o�;ѓF�V���&�K�5!o�d�����\����I���#�w�<��>�p�=�ހ�j1�W x�������4���\]\���hy��&��i�G7�o_����̀ʺ�t��ة����ـ�2���e
s�荞cT_B#�+p�"�F�1��Y��S2��G	_!�{�A�Հ={Gf��E�:S�}�R�<��ȇ�\�;>]+��cp��;�@^z����?,V�a6��u�a����r�	n5 @���|����k_[�'v0�R2�q��$m����3�P�v��;-��2P�s�7��*�e-�H��%��
o�Q'{�O����a�2h2�va���2��K-;�&�]Z���b[e��*	�<�$�OI�G���ھ;���=V�As�K��;�4�yK]�s�e�Vo���S��B�P0�R�^Jq�����p��*\�E�=���Y�+��R��R���J����Yl���^�R@��c�*��|��Y�;*%/9�>�H���{�"��z�墺~#��*4���J@�n�27�X�zP=J����[_��1&�E���Ly�I���`vK����y�w�LǀN2zg���e`��_�̴�X���� �H�8Ȉ�K����xZ���Ĉ0��l��E;����q�$<>7a�شB��`'���"=��[�"���v�����7:�~p,'6gP���x:�~Du�UI1����U��w��I��[8({>,n#v��}�۲�O6���'���=>y�H�Vc��}^:�~þI�>�Ҭ���I�X�s��$i�C�]Wk�'}��&�fA*X���C�j�Vu������Y�W�v�h9�Ui���.{�>�HYֹ�ZܤiM�y:2�ڋL�t	�&p���%Cj��R���c=�>_	�$�������XN�ɝ���-B���B�%^s�(tϷ}^��~"O��{��;���!I�f���Y���/8���"�d���nAǑ��s������΅�x�]����V6;o6>��7�ܤs�	�W���)\_�%��>3�|rW|�8z&&�%N3@9�u+�}w�9��6p/�a�%$0�e:�IjLEv��bй� �"d։����RsS��ՠ���!ɬ4��}�C䗑�Y5]��i��y�Z�s���f����xg�Бߧ�.B�;��Le7&�:"!
ň��GW�>��wc�4H�	M�;a��,�t��1ˑ 5E�U7a�'l�`,��"*H���wïY½�Bû��6�����Mc?hrPG��zc�A5p	X</���5�d��6F�E�~�n)z9�8Zi�_�^5�YY&���o���p�]]��u�1Z=��iy\g���8��}c�M��3��1�W�X�=�Ǚg��O��)��.�R��	�^x*���p|�Hp�@�9�0YTy�C����M�\��~i ��ƪJTu{��_����
%Z��gn�6x�8ye;<?H�Zqe`�
�M�U�$_ꅓ�PR�Ce>�Ow�2\�!��z�Q�L,���5�Ϊ���1�J8Wcǜo}����;��l���5��jߵ�Tͷ3�|��
?
�.k?��t�X�X�����Q�+���sB�ls�Q/q�H.xQ�k螙�*�ˌ����26�b,�>(xݺ�Xb�v��wrl�����iđIț�}�)� �l(K�h����y-;���Eu��b\Vz��3Ij\Xj��d�F�!K�^!�#T��X�����&��M�)��MǊ,�u�_�Y�|�1��S�n���Ź,%S#��SK7�`�D��It0B���J"�J�u}]veX*� ��䡈�K�;���n��~�7��	�N���n��=}��E�S��b!%�a�\�9���l9�Lە#�S� ��)RnzB~�Z�I/��������g����oyV�]Qh+�۷�}�<�z���1O�����1-��3$!b�h�b�t<8�Pt�	�jH��v�M[G�6:���n<�q�	���n���=R�n1�Vh:��߷Xi���⇣8��rW��W>�n��j!�h��x�����_H�9�f_b  wq�'sz*ފ ׊���B{=DUuss�n]���\ӷ��W�Fd�J8I��l}��O�]��VeRVi�����*i+��nF��3B��Н�uoDv�!w,��<:I�̈��c8͜G"e��xkBX�Rכ�������2�Q{�i��,����@4����'̝2�<����	ր�/�]����|@%�G?X��<�/k�Ab�CԗH �:��"+����Esh6 �(��I#z�{���b��Θ�'O�Y�x�b�����V�O����Ki\=�ʌ��C5�o�m���)����Д�ƙMat���>���v����;����}��c��C.�Mm�ҏ*�{�!����\��&bٰ���b*>�%{ב���o�1/�F�)4�B������j8�Rӭ!����$c^����A�a�[9V3]nn���+�;8�Cj޻�]Q�(������0:EJ;�Y/��J"���/�� 5-�?k���W �X=�R�:��/|�Q��V�8����A�8�������%���Ä���'�j�����?��li}��7Wc�@^��9�
%��B�ubNO���T�Z�Z5H ���g������� ����	r�AW	%?�1���AtP����!�lF6�o��M�c@g����{��I�|!�#��`�ٖ��C��L	0Wy0�L�G�N������V7�p�{-yKV�&�s�U�c��
��KʫL��]��ܜ�@;r��g��Y� X���R��Q>�/T��~[��
b�DV_!����s�e}�W���Nx|�{�'��գTDƧ�hq�����2��j�U����)s����f~G3�Di �o���o(">kG�`���P�'C�ξ��|;r�ƥl>U��[/e��`h1]oF��׌l�����L��8,"��p��z��Ze���$~��t�E��WtXΏ�r}�v��d�]3�Rl���Ο4O���t��x��ē�}�3	�<([���Bx���MU�{5��ck9��LY����#-E,�̗R�#!���Eole�>;��V;��u���y������P�"����NPQ'�i=(j-� X�����������Y��HdX(o�W��A9�R��i��@m�#ms���D5��V�1澖����h�I&svG�!��dNc����K+�m��bD�C:��R��R��e��-7f���ʽ~l����ѽXL-�X���Z9���P��#y0�j�T]��)Sk5�gŌw�k�Au�K�4Z����?�g�/����d���7�2s�ȶ#h됕��;�A����x\-C=�>FJ�Eڌ⮸�8��mBQ6�IK�"�*�pX�iQ�ʰg������B5���Ԣ�E�����	r�����,y>�I�(��S���x�1�E�X�+RGc�g��0�Ct���n�v,K�Y�;.������-��Yu b_.�m0+��#3>�l���X�&�P�/���.��.Ӑ)�Y��Et���]]~K�@�c]�͌��+PC(V��������e�ҸV�a���0�A���1�y��?�o���Q��<���A��{���J9��vu+��/z�I�uЯcN�V��b�@w5>�3$�y#6ǈ�\ =ΟH"���60/�!��e��`�w��m��m+c˸�I�7}��?F�w[�������4����=�mr������o�mW9�2ڗ/2,��������9�=�?(9�>r���Z]����ADX�A�p'c�q�#S!7ۉ��MN�  ��IyF��$a~G���R�q�%T���b�s(ܔfǨ��_&t>�m� ����OB.�N��9��`�vW/�
*�o~H��rpUl99%�+`[y0��)5��0�]��a���]������A/�7��߁��p���z|��S�����qi���
yI�H.N_ώɦ&��}�2el=��I�ִH`J�z�76v���".�[��exL�r{UE�s���U���ǜ���"�%�(d�3Q�"7�)�W-_�ژ�R���¬%�Ln\�Xy��R��qJz'���EIw���-�{��JS���)�>C������|��ոSC8���I��,�c�+�7�Y����RJT3�؋[U�H~���:nFY�Mq��jy��o��ߛ^���wY7�K��P%���l���6��9ݵ�u�}�_��`Mh2o����E�����q�=�%�S��ϱTM�@���J���$$e�bg���e��+�^�����`��7p�KY\�����7�]��8�<�
��qrm_��?���Z\(�� j��A�I܌�Y�6[�ɻNk~�������Z��xWX�9�=��{'sv�/U�Gx�[L�j�J�|h]/�*!��5y��%��n��_9*_�[		qN${����[����<C���Ӈ�6�T��Ǎ�`5C'��*��dx��/�ȫ��H{�����E�P���qA�����U����z5f'm��k��Bp�F�����]�s`���x���ǓB����U���T�g���k�
� y�w��Als2퍧��!�_�����ƹk��J#����+MD���ERrSɯ2o-k%ԬV#� �P��&&�\@_���G0��^��'�W�'�m�;�S>/2��2p4��`�@���2f��X�b��d���Dc��*N8�� �cBg��\�T쮘�6��;�7�,��+�VȂdܒ��EbZ�Ϭ��[0Nx���[ yl�]b��O,���5�2=�t������mE��\�r���1�pA����D���Zo�5� Ha�V(�ˠ�)�^α��n�W�������/��v�����Pz.&��@;���J�)^��F캇�[^�����Fo��U�#�\���Ƕ*ZkwW��Uz�[�N}-i���f1{��'Yjw�!���;��j��-�j�'� �hv���}\�v���&���f�i�P��S�n��
�&�]�]ꨣT(�N�g	كJٚc;G�Fܠ��9o�gHD���R�%8�I3JKmw�j�#p�b�YF+���iyJ�QCV6/i�-�W`�P�z4i�#ݵ/��ɉ�4/�N�^��U|�4\'\��I��G��6D�7Z~	�W�s�7�����Y�õ��j�4r�P���z�(m���r._�}�i[u%���|~P�Dh )uΏS%\�2����k��]��|��32�D>< ��d�Ɗ�t#�U5	dB�b�,�TCt�xhѐ�_U_�D*���$8o���lD;����԰�2�ւa9�f��L�e���mQ���)Ρ�_�*�i� H{y�Ϩ}�58�Lr7���q>�K�O�:{��B���و�5藷�7��{����FǮI�YS��5C'qذ�f��l�&��7nd\Z�Z��Ak�̐�,Zb��}3�i���~Rd�X��ȼY��ZZu�e!�� Kǀ� � ]"���{���(�z[�I2ѧa}k*�]�G�$a�WB�aP�'�=I6�?�p�>yI��XSBK>B�2��8�G�QA��M`o�� �(n����;���D�⽗�O�Mq�p���?)6J\m�M�=��p-�G�e��
�i��� oYg�O����X����}\c5�c�@��$�E7��$���ӑܑ�G��;IЬ\��v~����Y�4,��לǻi{)����O�@N��ɋh�T��5�P�%���wkfe�"�D�Y�O̮��~#�p�m58BN~��S<�.L����(	��fR�����O�F6g�(�R6p�@���ᏏGIJ.j�Zf:�'�߻-�_�iS�k���$�q�8�(߃`�J44h<Q��S{(������a�&{x���*�����v>�=��7D`�e��q{�xXie,Q�xq`�T~�i��š'�1�⌕"J~~V���Wޠ�A�;^�}FN�&^ѳX�s�1�O�)��쳣D��RN���#�pȲ�	� ����m���-)��+M��1'�y�����8�7&�é�񁫔=&Ou����d���k j8�B]� `� y������$\be�P}W��*[IR$#���=��;�N�F�D�JX�;'��=)��qAdE��o�U��
�UR�R!i2�o1����C����?^���g�#�@.f#��B�C/'�1eS�SG�N[����z��2cn�"���\���I�>�7@h�}�A�_|����X�+�ʒ^*���蜶r��a�O�B�����¶�M����U�v�w���g�Zx�������0u+�>�Z@Ϛ�
^'�9�~��'w�yZ���6R�[ӯ��Ew��>I����i�h�A���:ҽ�5�� lvo�{�z��d�`��3��-���5v�z�<���Ț&�8�?=�#�ә<"�9�b�����-"2Lۄ��3��m`W%��
�I���l0)t�ԫ��i�LfI7�F��J[�YVD�v��o�w0�>%��<*���zC�!�3Pv�п���؆j�,D��Qe m3�H�]
*\�d���D��nHX�ǅ�I�1���#+r��� <�h@+)pH��:��_s�}{�qD�|B�k�S�0.�.p~z9�P�����]�)�$Q���g�'���g��!<q^���=Y�L���|Mx`��k�l�	��v�%�QL��?h�ݍ{��~˸�`7r$壻oLR�IK;[�lF؝���Hb��36L�U���ٜ_0�PIw�ZS�̽-��}�:���mϤ5D�Ή��ę�l'�)ɛr�,笿|� �r1j"ɀ��;/��䩻(�$Y�J�P�9���#��ADBq��9P���hp�:>�#a&m�ݶ�8�\xv�~�r��8����G��T��À������WuX	�����zR�Ι��M�2&����%d��"���ط���hd�|[�� ���;�Z�nB�8� m���I�sb�/�5�\��q��FA'X�QG�0X:�6�j�\��qˬb�o��ːWH'ř��R����/���H��%{����(��Mԣl�ѵZv���%�=o���]�4�!�/��"�܂�-�Q��k[>��q�ɹ%.T=��������S��?�?��֣t�i5;c���g���T��zl��T�F��1$
���С�4�Pk�fC��`㬍[��^֜mǧ�q�Cyݾ���Au��4G��_��<N����z�˴�@.��}o(���۱
��,-��.�l�5���	��t�1�(���A'�j3�^Bq��QQ�4���	L-CZ�(o9�B��_*Qe18[�s3��i1�Xxh���ʖ�dG��3I��FQ���+im):�7T/(x�bR��<�PBb��A�s�$2M��Ҵ�][��)1�ivu�S�=o����KX���2@ր�X�D�j[�l������ȍ�p��(�T��[��l*j�4Ȫ3�j��Eq�q���U"�Wf���̤�׉]���x�;Rʝ������m���Ng��Xz�����6�~�H�w�?ҝ�%ܲ
�/�K�H�k�>QW9Z����PR��I3b��+�	�6��A�����Q?�M���� �:��Y�e)̷7G�*�/�̪�[��A�a�Z
��-��g��P�* m�l��/�"�f��8��?D���M�4����Q ��~��\e�{�e��AQ�}7,��j4��]���y������-�ڲ�ќ��i�rb��v�ʹ����w�f��.�|����MoC��UmAb/��_p�	Q����kc�eB	ޙJ��+��(/�x��v����P蘻v��w���:�	{q�B� ���fN�V��)�G�
\7 �����+�H'<�;���j��Z?��i�S���Z@I�KJ�C�ˇ &�<p�\��+m��Z#�M���k�Ք�&w�f��-n��������&$��ؚ��ƾ�6Q��e��sw��D�