��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����Y_��F��tw�p�^�=�����DW!of�.��"�"V�8��Ua}W#R�M�-Q�xq��ų�����#k_Q��?���B8I��c��l��{ͪNȽ�D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����~�Yp�����ݏG��@"�/�<��MI1|l �V�Ԕ�<�g���Y�L��]\.��{M0>��g�@����F�^]��p�)�L ���[z����;�6o�}�lb H����l���m���#SrRkyx����M��|9�
gֺ�(z�k� ���|Ok/���ԱJ���>�kP7�{X��A�M8�����;�踐ኜ�=u��!��r���Sl���w��s4���7�[���4��y��4YE�e�LmQS�ʞ��=���^_�1�b�t�6��7�B��\(��R���.X�	�������í�P>��uhʍrgJu��x�Ӏc�YҴ�����@|t����_���<�r�ƲP'A07����~է��!�?(Ucov�^���_���l	����;��Ԩ�{Js%M�Q2X,Ζ��f�"�(˼��,�n����[���.=�}�_�qJ���7���#������s��>��=�G��iҳ3ZF0�w�{�d$D��Uv�������N�m[D{T	D� ��c�(z�(X\"���39�oe�ͩ�Y83;e1���(_�����C�$�4���F.��)-�T,��5����?̛��oX�Y��e��IM���3�
vB�U
�1l�}䍦�D�x�Ѻl*��;)��G;����	0�9��<�ѓS�wN�u��T#/����1"}�^��FE�X�x���Z�i8�Zǩ���o�V�7xL�T���*�����[M��:�G�U��aY�xI%�(��J%������������Oť��|;����+��V���=dmL���(#@�m2eQ]�#�,�^�LS������>b��i�{/�٫�ɨȖ(���-��\��&�*�h�ǌ��	gޝ��7��BDndv@��ų-JҞtK��z��)�3Ϣ�%>�I1�P�*�:��<�:j��*�9�Ol/�pqf^��E�=��@%���_�o�@E��=؈a������#�iU62۞�t�p�$~/q`(	�g�,�RˑV?o���2=���3ǿo*`Q���l W����BkCle��A{�+�ɏVs� �F��P��W���3�|���n�q�i]+��2�t�����'H�w¬A�
�]�]B��<�ȫ�@[��9�e5�Xgj=� �v���Aa����fJV$B�<�c�!�sP����_inE�S�I9,lx�Hi}3cB��Z,�˳�����2~q�[`v(^x�f!X�f��|�f$(�{���[],k���a��!��5y���x�*��xy��"<x{��p�US�Ա�r�<0<�)X�5 ������}��_0�@v���>�����A&��z8�I6�Ƕ��#�YT ��M�@�o`�?5N�Z\��0������R6����^S�Au�%���됙4��`",�/R�X�8`.3*)�{��ܵ����p(��"�2��Y;�$�ϛs�A`��\�z�X��.��0���T�]el޾�TX����As:��P�sb��M��*ԧ�J���	S�E�ɼo/����T�u;2?����οl<.MiU28���,[MM�:�%֟l.f5o
���p�u�%WIu��w ��.���{�dhY��u�鎴`^��͙>I���xB!�*l۫hbi��}��l$�ÿ'1L@��1�/���>pbF�UU ��w�l�KvV�M�/��Eb�S�`H��z>0�Vq��TU�m�,ظ��y<X&*��aZ��0�ԎB_���G^���d�͡c�@��7��G�߲߇q�%	�S�����8��M|اB���VZ-��q��+)�<��o��g��@��r�����⟩J�1�gҀޢxr��\���B޷1�P�ȓb|�L�V[ݹ0�p�������
�z��ŏH�&,���%,XklgMC�
UJγ�W?���S<]�#�;�CkL]��S�~H18$U`�x|J�Fۯ���%~�UY����!˜����u��?��A�Ū.^g鴷�a�&�b"��Bаw�yL�;4��GA�b�GJbE����������^��(��5��Tu�Hs���▋�Wd�b�(�f����2\� ��sW��Dva,��d&Ʉ������t��]�z��(����ȭ�pv�3Z)n��ԕ E���HM���Ό�iA� V�f�6�cK_=���t�Z�R��U<������Q��|͞N��m��]C�*xI�6��_P;��z4�5O��S��Q�����H��+�����ҳ�T�����o(�l'��9Ҟ(W����(J�Hҷ���i>��M�X�� ��|��gܳ�['UB5	�C$���1 /�2�E�B/�%z!�)O�ȌM�~�xo�b�aֆ��#�D��xt�N��S�$s��j�
)�t�_L�q'��>�X�,
�a�=4S�Dl!������/� �������P��E2��?��޼���ɝ��.)XWߤ0u��/x5��w�7�����5�)�&�`��g�9�U�]�N��kQ�µ���r���e��R�_�E4h�9��;�%7K6� t����Xpۏr �8���8"@"���I�~P[Y�tܤҞ�������kopQD����u�"|��U������@T�D2���z�����6��qZ���}Eݭ��8yt��1�e�;�@���`�DɤĞ�q��ҿrQF�W�
�|o�-��$�x	/zQqhF�up���-vi~j�j���L���:p$Չx/�|��i���r�EW���M�qN\�Թc��$i�3�#}ɗsW븭c�T��#hJ��s����|�"���ֽ�t���g��k��N�Z�-5fO<6* Ŀ��3��Q|�cy.ښ
�	��o�і�m�Y�B��ހ����{�z줜�e6�~W�����iyfx<��/�V`1-,CP����هE����=�u�_?-��g�5g�����n�$�Q�#����p���bd&��eq����cB���g���v�V--���W9#��[�����/�^�a�%�]�Q�ݲ�5���X"�r���K}N?�I1����գ��� R�O�q�%���id�@��I.��Y ]��v֙=^\�śÒc�����+���kn�hGrpٝVΊ/5Zȣ��P* 4=�1l&��x���:z�:�.���d�-=���fR�h����c�%�%h���'X�1�|�{^o$����9@�7����m�-������<# �KO���]���p�J ['�2��.��M��.�<�"N!��Z�F���bD�f[���;��"fimvb�wA�
O*��Sټ��lW�,N)��D*�n��S~�z@�ăq9��(L����ܬ�l��_y8�2���M�'�o�a��J<7W+=��0��+�F�C�T��0U�[��CE[«�#���f�����x��g6|��TP�,ga�v���@>��ؙ�칞�ȟ�/*z�v�8)ߊ�C`�i�{\�M�n,q|ou
߼J�x����2f9�)�[U�zz�݈q��EMNR�s��K�e
���U#�׃Q#�@�o\~Ć�����˝ѓ9����!Lb�m�����'�O�N��wy�~�Bt2́��i�,͐�4x"j��3��@ �t�mLp�=����90=q��'�B �޼�|�J���v��d��"0��s��#�]��y���8]h����B!y9��i�&��Z�B���ٮJBR1�Β��I��0)��s�ɩ��ù8���hkMb)6�4�����|�hS|!�;D?��I/	�Z�% ��'\u�W=�7��v����"n���y�LPd�tRr�D�`�&�����+9`�y�?K�a�K����AWR��J��I6��7hS�&C�Hޢ�߃�Am>�O>h�[�%�������Nᅒh�󋎩�K�a�K��[�N�
E~��M �vݒχi�!r<�����|�lo4��h��S�@��'
p��N<er����M}�u�K���JuƝuJe��.w� ��:l��u�����l�J��2�!���
θ�Vc��[Lvf��r��6��"#�D+I�ӬDj2�:zfp��E Υ��8r������e�PN"ۥ�H�*�[�����|�̽hR��?wTE�T5*9�_���'p��i�VҢ~"�~�;s������J.M`��7��.�V���R�؞�M��V5k·b=�c��ΰ����>b)R�^1�)ʉXn�l10�Fm\u���}(]�+��ߦ�����B/d�9�q�{D��&9g""C&]d�)����l�*��?uCҞ��
���d��)�+rE�Q,�|�������u�/�l���ޗ<�aj1!A�f6�ѧ��u	� E�;������������}�^,�0��$]��u��hj�B��6&cN~kC(�h�h��ڒAR��v���m�5�)�������Y��b���o%M����X>ۤ��ڑ+�����x�n�3*e��;��b�*��P*x�b\>rn_Nd8�>��qLW�,�N)��KZ ��o5)�L��v����	���і�Ƃ\O]{y%a��F�]-Hu�o&u���mtK�������S:����t�t��(�c����|�eq���*Q�nߓ������:Vȥ�3V�:kⶻ~��n+<Ii�䯏$�`�m�fwbWL0
�G"��N���s=_�?��0�`؆�܁���gG+4���.�xk�m\l��V�w�f�c���7����Q��om�����Y̢�$�$�TO�~���w���[�n?ů:/���N�W|eHa<0YMף]�(돧Ȋ����y7���*��L�c�_T�Z�o�t̎gy3�XK��t,�Q�!��J�nd�	����D5��p�f6�
�2��c��}SO%0s�oB�i}b��l����&�*�S����$�=�$y�@�P����AV�.�3�Eer}]3]`�9�Ȅ)� �����-���)�	�|��Q��	2�\�)��r���]�cS�z�n����TF��,>�y���M�@�EV�Eq��=y���P>�^-R*|q����eF�?�M%�m1w���@���<��?g�9T8*�f�.��VY��6Z�u�#�t��f-!>R� ޚ��%9��Eៜ��xڕ���N�I�˝f{�(l���[��B��KR��P�g{�ߨȏ�\h�Dn�À5k�\_�+�����c�k��ވ�G�t:M|�ߚE�G�lb��snI�zw��d��L��ު�k�֭�Ͱ��R��+���c�ۑq����k�z*�5���?RI1�r���S븥�S�u�aJOԲnò�#�����-���s����'�5}�����,��^k��y+���S�}�`�}�y"�rD[Y�Z��[(n1�P����w��a��H�#�bm; ��K�&=0�P�Y��5l�2�5%\����ʹ�n��{Kx&D�� ~�x�@�L���U\�M!a�U�W���I�;+�a7��1�2W����a��f_��M�H���Qh..��Tm�Q\�ָL��j��|�8h���/��i��覻-m�=�B����'6�y�%`��?gan�`�Q�	�bq�3�x���Z絮�9�{�\�X��w�g���m
9��4-��&������������t�l\V~h���rV��\��CM�^o��O���.�u&Ƒ�d)�zOC�K]rW���������q�!��}�݂405U2�dE��»��:�i���nL�$_��s��kD�Jj��D,+{X= {�V�F��}l����9��u�=�I �c^؀�,� �U�ڬ#��W�hk}���G��s�>h*��bF,���U��xd^��~�j��ɱ5)^�w-���k�z6_úW���e��B�~�ض �|jd�����aBֻ\����Z� ���@�V��6�������>�[��lS���V��l���&麣��UÀ�prr�sZy��-��ה��= K���e����s9m�+E5f�6S�n�b�l9�~���eh��K-(r 0A3ڗ�MuA?X������!�;L	�JX���ޏ"�������ǌx��nM�ʯ�l�hF��u����$��YoȁvV���<�q���|͕�.�b�QpZhass�7�Op��y���@�|,��@Y�����Jq*K�1��+=L@�,���N-�<�e��P��H��8�_�$�}�U����`��0}�$f���J�*�r�<��H����e9#Z��/��nqk��d\|�h��xL��M���w�y����ֹ�D�z��HW��KM�gg�p���X�����y4��^�]$����D��B���$��Eůb9O��@�_�	��ݒ
�,�C7�=.��N�O��VԎ�.C��!_��RܷLD��Q��#�v%��,Z��5_�: C�+r�3dE (�C��]�G
�{��m�6mAkU�R���A�mD���c�w��b����WL%�N�*ɋ-���ș�.MxX*�R��U��߶�f�ZC�h|%�����־2��[3��X|�d�^A|��E!(�  ⢎��$��E�x�����q�ao��C1�ё�y\�G)�{8����m8/`pa)�R����
����_�29��(�S����h���̃��N�Us#!i! �9ɺ�j�V�fMT�&�ݶ��8%��AKԸcS-������*���=��N��$We4'��r�����!;��M�X����i�̢��M��L�QS	(_��/u����0ѫ83���&� �0|�Ԗ���0�ǡ�s��^GG�kǗ�e/���y<p{�����e^��j��Ē�#%W�~c��j�0�]��e�I���lw��=mz�֓�MGg�0��v;#fRX8��+�U�z��6���A�,��F�h�P��<��a1*���}cź1Α/�L�M��0e��"���rf�����ݛ)n����/��o���@�/շcg�z����w)P�7�^
�n�D^�F��򓇃�p��}�����^b>��k�Q��y�3���"pY�^��|zf��?�Ң�x�t�Q�p��iѯ�7��f���&��W��h,s!�\ ���8F�J�1T��Y��A��O�մW�F�`e$�]�@3?���H���n����B_k������W�#��5���"~\����d�Kܰ�~���>N����84�v-�mܞ���r%�۪�^Q�\��E�݂��S�h�g:4(�j�|�������
4�Ed~�@쨾rC0Ԕ���G����wz��?gb�ِE�1:�\�P�lfD���B���>r��1"Zc�:&�o��OˁM<��'�[R�.�C�N��.�/Ҧ��1��+п�97�al'֣��:�ZY����� �q������L�x��-��;�\A��T�^0N�e&%�j�p?4ucd�5���ӎ�5Ar����rMi7W���� �MCSϴ2�G˧,�y����V�� �R��p���!d�Z�J�p�7Oڤ��j�r�I��5��q�\z��0�&�5�Y���*(���ް�"�}�0)�Dی����T��1�W�����q�Lw�X���3���E��'|����OF�GO�1��,BQ�qڨd��4]@��We&��nm�R��B]��ő{D�W��� `y���N��z�0���\�%ez�t��U\L��"�!wl���i68�Pn�N��.�b[:
�A��D ����n�D8Me�ؖ[D��To�F#s����j��D��Ԝi�0ۀR���ט�Eenrf	m�� �(�k,��� �u\�Le��2��_{½��M�'ف��R^I{�|7D-����Tl[]TPam��G�ʧ��$'�$�tX�+cY4gZ��F��$X'��#%(�0y28��b ^l���ָe�Ÿ^�K�2�q�n}f����j�Ǳ�|46E��vi[�p��*#�����!��#F�2>��׊��F��>�s{.l@E�e[�Tm��S��N������yA�M� ��4�MF�d� f�pcR)��Qm8v�Ԏ���b���� ��9	f/6��B[9h������C������z��j�����/�x.q]�/��`0�A/�&����C��ƪ�.��M�E�*�,��v������v��'��Ƀ�Z��#[pNX8�G6S��S�ݥ�o�6Ci��tp���nS�&;_󴌛s��_��_9�P�����m���EV93U)�>����d`=)�P63?����}O��,o�n؍�"�z�jϡXA�b�u*�����}��ގ4zrB�\x]Kj�gf�F�[NͅO�1;�'�֧;�� ���6*RbuaA�w��ax���G� 0���Ű���!^隶f���D����a�``z�� #��e�$xZv��i~�Ð����h�9.gNC��I���
O��%����cp�.Vià`_�̓��%�4K�'�(�y�"N��d�_�|�#Ye��#tXZXE����)�%/�_����'�t����f�����d�i%ᗸ�fi��ٷ��08>|�����x�$a����x�:v���%�03X.;��CX�|�G�:�9$&�b����v�nM��}#�`�.���o�c�m-�ݳ$��]���=�*�r)C�Cl>����sB�"NEw����i�=��chU���*���K9[���wB� ��q(���0c�/*�(Y`?*�؜�� K�M�c����kQf<�'(�+�v ��R�I�n�c�i�&��lm����X!Z�8"�됯�03�C"uw���y~�9�m��K>���>(V}0"t�ۀ�3#��� �����ac �H�7�=��`�h9��G�r4��Ї@Z"����
��ApE*[����ߵy_򏶷�7�Β��+��)��]�œz-k�r�B����	�;��S����AX-�[�¶�&��^�L�S���~���qNk�٭��e��������C6�����׀�;\����*qC�ig/T�}���;9c9�v�F���e����*��&��+�a�Z�C��	�J�2~����]�6P�W���E臙"�Sx �pd��Ð�]�5Ŏ\��� ��䘻����f������hX��c��r*�Z$��5���<���ر{�I�cm�a��"��P݂ey%<����:t
�z�VQ��X��p=��[c�S�1jm�~jپ$��#X��y��mߗs�5�{��(_5 �&>Qi_.�ՙ=�KY%7��"I����6"�t��w�H0�^3�k󛔬�Ϗɤj�����x,���9��y�<`�L�EbW��9��y�U���T�9`�.�n[�7�6���u�`�	[�1�1������d��BnB�&��� X����<�������jRW��W��ٝ�7~Q����
x�,# ��z:���,���O�]Ʋ6��)wV�5��q`~u�]���Ԇ���D��G"����M��}�>"�\�<�ms���I����-%�j�v�jY�|XuU��8D�A��h;�l���K�]_ά��*�X���gh=9n���&����̴�p^:��1�5�e�u�\9zPj2��z���:X�L�{�n����^��'��?<���u��u�@C[cU�*�`��S�1H���b́��~ž0Z.w'�1b�h��A5q����������tf7�ێ&~ w��|�Ԥ����Q�u�L,KD+�*�y7�N<-92ܰC`��ǮH#�ٳW�s��8��L���G�h��	Ռ#4d6�WEkM�>t�4����Jz>��W�7��jp����ܬ?��j�)="R��7�7�2��q0;����	�J9*�6�-a������*l@�}�p���e;�b'�Υ�I�s��uG\�Rl��\tu��ңi��wXy�4δ�A5˗���H�|s�:�5.��߼n���CL���[�۷-Y��~���Q����raQ�!H�ihvr\"MD�*�ǥ8e��phvѺ�f^t�L�q������b$�ٸKT&[uvM[��vÜl�ٟ�!�G�|��IKɑ�>�c��쉒c��@�ӽX<dB���Rg��;��h���z(E�7p�$2C�X鳜�ۤqT֬� �u��q�{~ Y˒C��^K�&�Of�8*���ݰ�>R��/'�ʃ^w�^L&�N�ݧ�8 �m��l��У8�;%�aD.<�ے�\��؆#����-�d[��Ki�w����q�$����20n�,�ѬU���J��6�������r��kǦeҟ�������'������o����TG/P���|vb��n3�
�mpq�
B�Ph.u����d�`3Pϭ�l��urI@v�R6tx�Ͷ,��Q��Z�;�H��;�΅l)�5$��R�����Q@a������F�G:��-(��~��TRG @����������w�XBo��(��9�?}�$扐�& �����#��枥�#x�|�_�9�zK�5�>T�e�B����ޮ�X\�ڰ�����~����|��<�]5z��7,�[�Π%XW�sK���k��盵�y��R���26C��x��݈�v���6��¥o�e%��݉)�vL=KD\z�7�
�-k7�۵ռ��W����4��&Qr�GƔj��9�$�l�4Q�����Q�T��V��{�y;�-�ӄ����3lh��!�j.Cv$�n�=8��s顅�}�eн�-Ep>�,wH�^tM�4�d�Vn�g�8��u�*��uk�!�����_���V�����s!�3d!Q/��䔄�ã��c-��A�0�sa����{]����B  ��˼*R@(��?>*K���'��&�@�k�I06;�0h��م�R$����\2��C�݇�&�7CD&RۛUqk�j铩��|sD�#��.��7lc�Q_S)�kEEw���J��E�R���������AATO�&�	�v�(�{Ot-�,�(`�����/��by���:���T/_���Q�5�SQ�����3[�j����|�޵�� Xk��;�7!�S��@��Τ�Z�e�vJ�Pr�<�H�p��n�&W^,�7G�S�#:�\��\�����WO���q�42�p�N.�z���{9ɍ��r���í
wP���!��o킊�a4�jG:��ᦝk��RPD>��Q�~����r1���s0:0K@�g�V13:U��ڔ�}�PC���i���._�V�{�x�f�΢���^k�����'��Zz��]��ޡ[���m�q�ꏎ�o���P*K�1��yt�{��YO7qG��>	Oqjkr��\��Qٓ&�����v�nh����̎m��|�{b`RHN��s,v��:?e�(�V
��Y�HP-G��I���*
�C�:*xIHT�aD���Jw�m��b�2>p�YK��C�g�uI'��E7Ļ-7=����W���%���R�q��ܽ)��C]@����a���;�ek=|h��#k�`�}�ݣͫ�T�9�>_=�"�O����Z��`���LX�9�{N���U!�~���G��?���]�Q�;�rjO��OY���w����Ob����_�&ޗD/FS��ՠ+nlw�=���h���~��[i���qmHg��F>���k�9\x������Y�ν�]+i\�{>Di�6���p�������Ȣ��o4^:k��7�1�K/�[���e��ɤ�b?w@�;d��"ښ-��y�D����"�������Ϣ�H>PsM �sRs3{�s��26�3�&W�1����䤞�z�ʶ�L����S\x����]&�����ZY�>id��3���3�Q>?�!X���&w��|y�6 =���!8�n�L`/� �