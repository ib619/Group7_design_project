��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���d3�q	��9/�I�w`W?ދ�S"K7��5�,l��C���
@E=D��!
����荾Z�V�h��c,Dt��&�����]4w9K_9O�=l�uE�w����[R�\�zÚ�-J�$����åCj�[�
����T=���K���h�����,������#�z~��?�G���B�~֨1)��k��yq�$/ju�YA9��SX�{@��mWt������w�F��r���������O)�mC�&�����$��^_��|�����=������A���_"�s���50��-�ݡ��kVE~�cu��'Ah%�����v2ݲK:|�g���7/��=Q�u�~��qC���
qSa�a�n�m(�]�h-�FK�]�Z<��K�b�s��'�����C$Yכֿ��h|�[@lXJ�*Qm?�аR��(�v�vlr�j)ڦ��0p�s�bv��jy�-����(��N�vהS��Y�n)!��\|9��;#�o:�#��9|TWL��L2=�'���$ƫ���19�?�:H�A���T秧���,rJ$�p}�a�ڡ�rn#9���~�1e�[e���!������{�T�7���O�z�������쉎�<o�j��D�7��lS�ƃ���F�V�:¦?�,�:4I~P�o6����2
�ԫ�#��G롔�qH���'> x������>I�nN1.�yφ�V�ǹW�)��	�3���k��c�Rw�buRA�8����\��L+pȟ�U���R�z�]����X�`��.�2ָi�FeG��[>��V��cp��kɝܫ �\r6޽����8-h�\{����r�&?��e��gE�a�-�o��Ty,і65O$�H����i�������NҶ9ϕ�Ŝ�|~��	'^pڟ��K����B�w�o�g)��l)�L�'��|��<�zP��f��%"m�V�
�eR��I�3��%�`�Ss'�'4v���
�g޻�H2�~�)Gp<��.2������02a'�M�ԮNq%�$h�d��1x��zuק޵?ޗ�ρAt����i�����#��Һl0��S
!d���o@�9��g���=�)U��㕢o ͋�N,j3 1�*�bH�GH��^-[��B�>�G�l��uc'Xҳ�=<����Qs���ق)��!d�Ca�9��&r����JR�ff�D:�;!A���1�o�A�4L�������֡�L����d��0�9���B�x(�� ���d^�9O�
�񱺗�7*xȨkÈS����K;9@�_��3q�s�rc�P���^��*�V�zۦ�IR���L��c��q�/[LCZ���f!�N 6�c�������$j{gw�����	V�WL��xE��-����ͬ8Q�������>�.���U������h`Yj������/��6�슡~�&�����BaP3�ˀ���z�o�w%�s�[���q���u�T�5�ӹ�k$g��:���&"�C����6���UE�[OD�MD:��K�3��\��XL����Km���B(�έ��U	�Jܖ �C�~���4Yd^�CX���-G�ۤen����ϡ��6濡��n����U�����˼���"dV�w4B�M��4��%�i2��;�Ǆvzs��N�W��o���2��f�G��@#d[�[X�ug�|~�����/p��iɘY�  �����i��x��t���̅��R���,���F�J?���P69�\�W3�!�fz�"�Sw��x��)�X��(�`����t��;0�E�>�̞�L:)�.�����6��>���u3kH��xW�ɡ�0�����8�V�%�4<+)K�ن��y��\��R2�yX9K���;������<Y�������F��ǟ�ݽ��y%��>"���CEK�V�}���i�,��F���~�}��NFw�N!�x�,��nJ_<����}��5���=o���m��]�-�E���6�2��m��A�l˙稤��^~��7H�'�{i)#�XN\+Aaa0����V[�����̩O��Ϡ\cV�&�NzF�Ś�/]����"��X�yFe��������cjo�Q��1�l���"-������p����C�;<�s�S�P�{v�����k���<�GJM/��^����1��^�����i��alJFf5���'�?��ŵ�ag��� KX���!��7�]������Id�����D�k���u��ćTK�	_�&Ȓ�7�ླ�����|���>o},@D�)�8��w��Lb�Q�|��?�!���+�S�~�Cͮ��n���@��v 4�:1i
�+cѿ�o���Co�onp3�t��L&%h8��.�2��o�}�-���A�e��	��y=� o��i��Z�t��C��I/�X\zo���	�<p��P�*)�+$ْ�Ͷ��Bj�)�
�×��I�7���u�Xg�)���{���k�T�T?���E�Vy36�U#GI�a��a�	&�|������~1�,�}������G�Q��Q%}�/Py�n�Y�k��C�����=A�s�!/C��+����sh+O�����_uQ���!FN�Zq��m�0G �KiI��	P
:���=y�L�8ܛ�Ng�~_Mh��.��Kp&5:�vP��v�T�*��`�6��P�/G%����6�|t0k���d�b˨s0 �瘮�f�&�R����%"��q~\G���]�s��8���;�K5N�����j�j��.��]i����l��$�D����_��-)�l{�O��9�Z�)��|WV����d������<��� �6�F>�8�D	��ZF�C�J)�m��/2�����kq�S�%u�05��/�at����f�1��J
X�*A����K,������);��N��5�2�羠s��N�s�[O.�T�w<��}%Hء �l10���`1��D���J�{t��M����u��&��y-5w/T=*G8�f�Ǉ�O+M�jH�o�qh׏rp�.[����#,��KF�7�W�WG�{	�945�� �&O�6^����Ԫs�1���9I��l�2N��x����<_\